VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO wrapped_asic_watch
  CLASS BLOCK ;
  FOREIGN wrapped_asic_watch ;
  ORIGIN 0.000 0.000 ;
  SIZE 220.000 BY 220.000 ;
  PIN active
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 71.710 0.000 72.270 4.000 ;
    END
  END active
  PIN io_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 153.420 4.000 154.620 ;
    END
  END io_in[0]
  PIN io_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 9.150 216.000 9.710 220.000 ;
    END
  END io_in[10]
  PIN io_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 216.000 201.020 220.000 202.220 ;
    END
  END io_in[11]
  PIN io_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 10.990 216.000 11.550 220.000 ;
    END
  END io_in[12]
  PIN io_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 80.910 216.000 81.470 220.000 ;
    END
  END io_in[13]
  PIN io_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 113.110 0.000 113.670 4.000 ;
    END
  END io_in[14]
  PIN io_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 90.110 216.000 90.670 220.000 ;
    END
  END io_in[15]
  PIN io_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 204.190 216.000 204.750 220.000 ;
    END
  END io_in[16]
  PIN io_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 67.110 0.000 67.670 4.000 ;
    END
  END io_in[17]
  PIN io_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 92.220 4.000 93.420 ;
    END
  END io_in[18]
  PIN io_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 216.000 196.940 220.000 198.140 ;
    END
  END io_in[19]
  PIN io_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 209.180 4.000 210.380 ;
    END
  END io_in[1]
  PIN io_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 48.710 0.000 49.270 4.000 ;
    END
  END io_in[20]
  PIN io_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 115.870 216.000 116.430 220.000 ;
    END
  END io_in[21]
  PIN io_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 103.910 0.000 104.470 4.000 ;
    END
  END io_in[22]
  PIN io_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 15.590 216.000 16.150 220.000 ;
    END
  END io_in[23]
  PIN io_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 216.000 25.580 220.000 26.780 ;
    END
  END io_in[24]
  PIN io_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 216.000 156.140 220.000 157.340 ;
    END
  END io_in[25]
  PIN io_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.790 0.000 209.350 4.000 ;
    END
  END io_in[26]
  PIN io_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 123.500 4.000 124.700 ;
    END
  END io_in[27]
  PIN io_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 64.350 216.000 64.910 220.000 ;
    END
  END io_in[28]
  PIN io_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 24.790 0.000 25.350 4.000 ;
    END
  END io_in[29]
  PIN io_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 139.820 4.000 141.020 ;
    END
  END io_in[2]
  PIN io_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 29.660 4.000 30.860 ;
    END
  END io_in[30]
  PIN io_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 129.670 216.000 130.230 220.000 ;
    END
  END io_in[31]
  PIN io_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 138.870 0.000 139.430 4.000 ;
    END
  END io_in[32]
  PIN io_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 216.000 186.060 220.000 187.260 ;
    END
  END io_in[33]
  PIN io_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 133.020 4.000 134.220 ;
    END
  END io_in[34]
  PIN io_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 9.150 0.000 9.710 4.000 ;
    END
  END io_in[35]
  PIN io_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 88.140 4.000 89.340 ;
    END
  END io_in[36]
  PIN io_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 216.000 55.500 220.000 56.700 ;
    END
  END io_in[37]
  PIN io_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 59.750 216.000 60.310 220.000 ;
    END
  END io_in[3]
  PIN io_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 20.190 216.000 20.750 220.000 ;
    END
  END io_in[4]
  PIN io_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 83.670 0.000 84.230 4.000 ;
    END
  END io_in[5]
  PIN io_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 164.630 216.000 165.190 220.000 ;
    END
  END io_in[6]
  PIN io_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 143.470 216.000 144.030 220.000 ;
    END
  END io_in[7]
  PIN io_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 57.910 216.000 58.470 220.000 ;
    END
  END io_in[8]
  PIN io_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 216.000 214.620 220.000 215.820 ;
    END
  END io_in[9]
  PIN io_oeb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 190.390 216.000 190.950 220.000 ;
    END
  END io_oeb[0]
  PIN io_oeb[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 116.700 4.000 117.900 ;
    END
  END io_oeb[10]
  PIN io_oeb[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 173.830 216.000 174.390 220.000 ;
    END
  END io_oeb[11]
  PIN io_oeb[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 216.000 162.940 220.000 164.140 ;
    END
  END io_oeb[12]
  PIN io_oeb[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 171.100 4.000 172.300 ;
    END
  END io_oeb[13]
  PIN io_oeb[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 216.000 97.660 220.000 98.860 ;
    END
  END io_oeb[14]
  PIN io_oeb[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 22.950 0.000 23.510 4.000 ;
    END
  END io_oeb[15]
  PIN io_oeb[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 194.990 0.000 195.550 4.000 ;
    END
  END io_oeb[16]
  PIN io_oeb[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 48.710 216.000 49.270 220.000 ;
    END
  END io_oeb[17]
  PIN io_oeb[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 119.420 4.000 120.620 ;
    END
  END io_oeb[18]
  PIN io_oeb[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 216.000 48.700 220.000 49.900 ;
    END
  END io_oeb[19]
  PIN io_oeb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 43.260 4.000 44.460 ;
    END
  END io_oeb[1]
  PIN io_oeb[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 106.670 216.000 107.230 220.000 ;
    END
  END io_oeb[20]
  PIN io_oeb[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 82.750 216.000 83.310 220.000 ;
    END
  END io_oeb[21]
  PIN io_oeb[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 85.510 0.000 86.070 4.000 ;
    END
  END io_oeb[22]
  PIN io_oeb[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2.460 4.000 3.660 ;
    END
  END io_oeb[23]
  PIN io_oeb[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 62.510 0.000 63.070 4.000 ;
    END
  END io_oeb[24]
  PIN io_oeb[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 185.790 0.000 186.350 4.000 ;
    END
  END io_oeb[25]
  PIN io_oeb[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 137.100 4.000 138.300 ;
    END
  END io_oeb[26]
  PIN io_oeb[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 216.000 118.060 220.000 119.260 ;
    END
  END io_oeb[27]
  PIN io_oeb[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 213.390 0.000 213.950 4.000 ;
    END
  END io_oeb[28]
  PIN io_oeb[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 164.630 0.000 165.190 4.000 ;
    END
  END io_oeb[29]
  PIN io_oeb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 65.020 4.000 66.220 ;
    END
  END io_oeb[2]
  PIN io_oeb[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 216.000 131.660 220.000 132.860 ;
    END
  END io_oeb[30]
  PIN io_oeb[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 50.550 0.000 51.110 4.000 ;
    END
  END io_oeb[31]
  PIN io_oeb[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 85.510 216.000 86.070 220.000 ;
    END
  END io_oeb[32]
  PIN io_oeb[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 187.630 216.000 188.190 220.000 ;
    END
  END io_oeb[33]
  PIN io_oeb[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 216.000 135.740 220.000 136.940 ;
    END
  END io_oeb[34]
  PIN io_oeb[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 102.070 0.000 102.630 4.000 ;
    END
  END io_oeb[35]
  PIN io_oeb[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 216.150 0.000 216.710 4.000 ;
    END
  END io_oeb[36]
  PIN io_oeb[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 44.110 0.000 44.670 4.000 ;
    END
  END io_oeb[37]
  PIN io_oeb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 216.000 45.980 220.000 47.180 ;
    END
  END io_oeb[3]
  PIN io_oeb[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 103.910 216.000 104.470 220.000 ;
    END
  END io_oeb[4]
  PIN io_oeb[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 184.700 4.000 185.900 ;
    END
  END io_oeb[5]
  PIN io_oeb[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 16.060 4.000 17.260 ;
    END
  END io_oeb[6]
  PIN io_oeb[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 111.270 216.000 111.830 220.000 ;
    END
  END io_oeb[7]
  PIN io_oeb[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 202.350 0.000 202.910 4.000 ;
    END
  END io_oeb[8]
  PIN io_oeb[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 216.000 107.180 220.000 108.380 ;
    END
  END io_oeb[9]
  PIN io_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 57.910 0.000 58.470 4.000 ;
    END
  END io_out[0]
  PIN io_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 9.260 4.000 10.460 ;
    END
  END io_out[10]
  PIN io_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 67.110 216.000 67.670 220.000 ;
    END
  END io_out[11]
  PIN io_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 167.390 0.000 167.950 4.000 ;
    END
  END io_out[12]
  PIN io_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 211.900 4.000 213.100 ;
    END
  END io_out[13]
  PIN io_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 216.000 113.980 220.000 115.180 ;
    END
  END io_out[14]
  PIN io_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 216.000 217.340 220.000 218.540 ;
    END
  END io_out[15]
  PIN io_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 108.510 216.000 109.070 220.000 ;
    END
  END io_out[16]
  PIN io_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 216.000 158.860 220.000 160.060 ;
    END
  END io_out[17]
  PIN io_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 176.590 216.000 177.150 220.000 ;
    END
  END io_out[18]
  PIN io_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 213.390 216.000 213.950 220.000 ;
    END
  END io_out[19]
  PIN io_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 71.710 216.000 72.270 220.000 ;
    END
  END io_out[1]
  PIN io_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 216.000 39.180 220.000 40.380 ;
    END
  END io_out[20]
  PIN io_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 152.670 216.000 153.230 220.000 ;
    END
  END io_out[21]
  PIN io_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 216.150 216.000 216.710 220.000 ;
    END
  END io_out[22]
  PIN io_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 112.620 4.000 113.820 ;
    END
  END io_out[23]
  PIN io_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 190.390 0.000 190.950 4.000 ;
    END
  END io_out[24]
  PIN io_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 216.000 41.900 220.000 43.100 ;
    END
  END io_out[25]
  PIN io_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 152.670 0.000 153.230 4.000 ;
    END
  END io_out[26]
  PIN io_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 38.590 216.000 39.150 220.000 ;
    END
  END io_out[27]
  PIN io_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 134.270 0.000 134.830 4.000 ;
    END
  END io_out[28]
  PIN io_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 15.590 0.000 16.150 4.000 ;
    END
  END io_out[29]
  PIN io_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 18.350 216.000 18.910 220.000 ;
    END
  END io_out[2]
  PIN io_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 216.000 77.260 220.000 78.460 ;
    END
  END io_out[30]
  PIN io_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 45.950 0.000 46.510 4.000 ;
    END
  END io_out[31]
  PIN io_out[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 178.430 0.000 178.990 4.000 ;
    END
  END io_out[32]
  PIN io_out[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 143.900 4.000 145.100 ;
    END
  END io_out[33]
  PIN io_out[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 215.980 4.000 217.180 ;
    END
  END io_out[34]
  PIN io_out[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 127.830 216.000 128.390 220.000 ;
    END
  END io_out[35]
  PIN io_out[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 160.030 216.000 160.590 220.000 ;
    END
  END io_out[36]
  PIN io_out[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 33.990 0.000 34.550 4.000 ;
    END
  END io_out[37]
  PIN io_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 216.000 179.260 220.000 180.460 ;
    END
  END io_out[3]
  PIN io_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 132.430 216.000 132.990 220.000 ;
    END
  END io_out[4]
  PIN io_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 129.670 0.000 130.230 4.000 ;
    END
  END io_out[5]
  PIN io_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 146.230 0.000 146.790 4.000 ;
    END
  END io_out[6]
  PIN io_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 80.910 0.000 81.470 4.000 ;
    END
  END io_out[7]
  PIN io_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 148.070 216.000 148.630 220.000 ;
    END
  END io_out[8]
  PIN io_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 216.000 120.780 220.000 121.980 ;
    END
  END io_out[9]
  PIN la1_data_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 216.000 28.300 220.000 29.500 ;
    END
  END la1_data_in[0]
  PIN la1_data_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 76.310 216.000 76.870 220.000 ;
    END
  END la1_data_in[10]
  PIN la1_data_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 24.790 216.000 25.350 220.000 ;
    END
  END la1_data_in[11]
  PIN la1_data_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 36.750 216.000 37.310 220.000 ;
    END
  END la1_data_in[12]
  PIN la1_data_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 167.020 4.000 168.220 ;
    END
  END la1_data_in[13]
  PIN la1_data_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 85.420 4.000 86.620 ;
    END
  END la1_data_in[14]
  PIN la1_data_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 58.220 4.000 59.420 ;
    END
  END la1_data_in[15]
  PIN la1_data_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 33.740 4.000 34.940 ;
    END
  END la1_data_in[16]
  PIN la1_data_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 204.190 0.000 204.750 4.000 ;
    END
  END la1_data_in[17]
  PIN la1_data_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 216.000 149.340 220.000 150.540 ;
    END
  END la1_data_in[18]
  PIN la1_data_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 10.990 0.000 11.550 4.000 ;
    END
  END la1_data_in[19]
  PIN la1_data_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 164.300 4.000 165.500 ;
    END
  END la1_data_in[1]
  PIN la1_data_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 73.550 0.000 74.110 4.000 ;
    END
  END la1_data_in[20]
  PIN la1_data_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.790 216.000 209.350 220.000 ;
    END
  END la1_data_in[21]
  PIN la1_data_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 88.270 216.000 88.830 220.000 ;
    END
  END la1_data_in[22]
  PIN la1_data_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 169.230 0.000 169.790 4.000 ;
    END
  END la1_data_in[23]
  PIN la1_data_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 68.950 216.000 69.510 220.000 ;
    END
  END la1_data_in[24]
  PIN la1_data_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 22.860 4.000 24.060 ;
    END
  END la1_data_in[25]
  PIN la1_data_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 216.000 62.300 220.000 63.500 ;
    END
  END la1_data_in[26]
  PIN la1_data_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 195.580 4.000 196.780 ;
    END
  END la1_data_in[27]
  PIN la1_data_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 216.000 207.820 220.000 209.020 ;
    END
  END la1_data_in[28]
  PIN la1_data_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1.790 216.000 2.350 220.000 ;
    END
  END la1_data_in[29]
  PIN la1_data_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 175.180 4.000 176.380 ;
    END
  END la1_data_in[2]
  PIN la1_data_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 150.830 0.000 151.390 4.000 ;
    END
  END la1_data_in[30]
  PIN la1_data_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 181.190 0.000 181.750 4.000 ;
    END
  END la1_data_in[31]
  PIN la1_data_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 216.000 104.460 220.000 105.660 ;
    END
  END la1_data_in[3]
  PIN la1_data_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 117.710 216.000 118.270 220.000 ;
    END
  END la1_data_in[4]
  PIN la1_data_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 211.550 0.000 212.110 4.000 ;
    END
  END la1_data_in[5]
  PIN la1_data_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 197.750 0.000 198.310 4.000 ;
    END
  END la1_data_in[6]
  PIN la1_data_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 120.470 216.000 121.030 220.000 ;
    END
  END la1_data_in[7]
  PIN la1_data_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 216.000 7.900 220.000 9.100 ;
    END
  END la1_data_in[8]
  PIN la1_data_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 36.460 4.000 37.660 ;
    END
  END la1_data_in[9]
  PIN la1_data_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 216.000 10.620 220.000 11.820 ;
    END
  END la1_data_out[0]
  PIN la1_data_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 191.500 4.000 192.700 ;
    END
  END la1_data_out[10]
  PIN la1_data_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 27.550 216.000 28.110 220.000 ;
    END
  END la1_data_out[11]
  PIN la1_data_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 81.340 4.000 82.540 ;
    END
  END la1_data_out[12]
  PIN la1_data_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 32.150 0.000 32.710 4.000 ;
    END
  END la1_data_out[13]
  PIN la1_data_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 115.870 0.000 116.430 4.000 ;
    END
  END la1_data_out[14]
  PIN la1_data_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 181.190 216.000 181.750 220.000 ;
    END
  END la1_data_out[15]
  PIN la1_data_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 92.870 216.000 93.430 220.000 ;
    END
  END la1_data_out[16]
  PIN la1_data_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 216.000 127.580 220.000 128.780 ;
    END
  END la1_data_out[17]
  PIN la1_data_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 50.060 4.000 51.260 ;
    END
  END la1_data_out[18]
  PIN la1_data_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 216.000 169.740 220.000 170.940 ;
    END
  END la1_data_out[19]
  PIN la1_data_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 113.110 216.000 113.670 220.000 ;
    END
  END la1_data_out[1]
  PIN la1_data_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 67.740 4.000 68.940 ;
    END
  END la1_data_out[20]
  PIN la1_data_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 32.150 216.000 32.710 220.000 ;
    END
  END la1_data_out[21]
  PIN la1_data_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 62.510 216.000 63.070 220.000 ;
    END
  END la1_data_out[22]
  PIN la1_data_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 202.380 4.000 203.580 ;
    END
  END la1_data_out[23]
  PIN la1_data_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 160.220 4.000 161.420 ;
    END
  END la1_data_out[24]
  PIN la1_data_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 216.000 111.260 220.000 112.460 ;
    END
  END la1_data_out[25]
  PIN la1_data_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 216.000 124.860 220.000 126.060 ;
    END
  END la1_data_out[26]
  PIN la1_data_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 198.300 4.000 199.500 ;
    END
  END la1_data_out[27]
  PIN la1_data_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 196.830 216.000 197.390 220.000 ;
    END
  END la1_data_out[28]
  PIN la1_data_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 216.000 84.060 220.000 85.260 ;
    END
  END la1_data_out[29]
  PIN la1_data_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 76.310 0.000 76.870 4.000 ;
    END
  END la1_data_out[2]
  PIN la1_data_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 13.750 216.000 14.310 220.000 ;
    END
  END la1_data_out[30]
  PIN la1_data_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 171.990 216.000 172.550 220.000 ;
    END
  END la1_data_out[31]
  PIN la1_data_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 94.940 4.000 96.140 ;
    END
  END la1_data_out[3]
  PIN la1_data_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 26.940 4.000 28.140 ;
    END
  END la1_data_out[4]
  PIN la1_data_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 79.070 0.000 79.630 4.000 ;
    END
  END la1_data_out[5]
  PIN la1_data_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 160.030 0.000 160.590 4.000 ;
    END
  END la1_data_out[6]
  PIN la1_data_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 216.000 142.540 220.000 143.740 ;
    END
  END la1_data_out[7]
  PIN la1_data_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 173.830 0.000 174.390 4.000 ;
    END
  END la1_data_out[8]
  PIN la1_data_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 101.740 4.000 102.940 ;
    END
  END la1_data_out[9]
  PIN la1_oenb[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 4.550 0.000 5.110 4.000 ;
    END
  END la1_oenb[0]
  PIN la1_oenb[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 29.390 0.000 29.950 4.000 ;
    END
  END la1_oenb[10]
  PIN la1_oenb[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 40.540 4.000 41.740 ;
    END
  END la1_oenb[11]
  PIN la1_oenb[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 134.270 216.000 134.830 220.000 ;
    END
  END la1_oenb[12]
  PIN la1_oenb[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 125.070 0.000 125.630 4.000 ;
    END
  END la1_oenb[13]
  PIN la1_oenb[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 59.750 0.000 60.310 4.000 ;
    END
  END la1_oenb[14]
  PIN la1_oenb[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 118.630 0.000 119.190 4.000 ;
    END
  END la1_oenb[15]
  PIN la1_oenb[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 216.000 21.500 220.000 22.700 ;
    END
  END la1_oenb[16]
  PIN la1_oenb[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 218.700 4.000 219.900 ;
    END
  END la1_oenb[17]
  PIN la1_oenb[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 123.230 0.000 123.790 4.000 ;
    END
  END la1_oenb[18]
  PIN la1_oenb[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 162.790 216.000 163.350 220.000 ;
    END
  END la1_oenb[19]
  PIN la1_oenb[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 158.190 0.000 158.750 4.000 ;
    END
  END la1_oenb[1]
  PIN la1_oenb[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 216.000 59.580 220.000 60.780 ;
    END
  END la1_oenb[20]
  PIN la1_oenb[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 217.990 216.000 218.550 220.000 ;
    END
  END la1_oenb[21]
  PIN la1_oenb[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 216.000 32.380 220.000 33.580 ;
    END
  END la1_oenb[22]
  PIN la1_oenb[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 157.500 4.000 158.700 ;
    END
  END la1_oenb[23]
  PIN la1_oenb[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 216.000 176.540 220.000 177.740 ;
    END
  END la1_oenb[24]
  PIN la1_oenb[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 176.590 0.000 177.150 4.000 ;
    END
  END la1_oenb[25]
  PIN la1_oenb[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 199.590 216.000 200.150 220.000 ;
    END
  END la1_oenb[26]
  PIN la1_oenb[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 148.070 0.000 148.630 4.000 ;
    END
  END la1_oenb[27]
  PIN la1_oenb[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 141.630 216.000 142.190 220.000 ;
    END
  END la1_oenb[28]
  PIN la1_oenb[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 20.190 0.000 20.750 4.000 ;
    END
  END la1_oenb[29]
  PIN la1_oenb[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 6.390 216.000 6.950 220.000 ;
    END
  END la1_oenb[2]
  PIN la1_oenb[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 90.110 0.000 90.670 4.000 ;
    END
  END la1_oenb[30]
  PIN la1_oenb[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 43.190 216.000 43.750 220.000 ;
    END
  END la1_oenb[31]
  PIN la1_oenb[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 41.350 0.000 41.910 4.000 ;
    END
  END la1_oenb[3]
  PIN la1_oenb[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 155.430 0.000 155.990 4.000 ;
    END
  END la1_oenb[4]
  PIN la1_oenb[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 146.230 216.000 146.790 220.000 ;
    END
  END la1_oenb[5]
  PIN la1_oenb[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 216.000 194.220 220.000 195.420 ;
    END
  END la1_oenb[6]
  PIN la1_oenb[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 78.150 216.000 78.710 220.000 ;
    END
  END la1_oenb[7]
  PIN la1_oenb[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 45.950 216.000 46.510 220.000 ;
    END
  END la1_oenb[8]
  PIN la1_oenb[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 150.830 216.000 151.390 220.000 ;
    END
  END la1_oenb[9]
  PIN vccd1
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 206.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 206.960 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 206.960 ;
    END
  END vssd1
  PIN wb_clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 192.230 0.000 192.790 4.000 ;
    END
  END wb_clk_i
  PIN wb_rst_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 123.230 216.000 123.790 220.000 ;
    END
  END wb_rst_i
  PIN wbs_ack_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 216.000 3.820 220.000 5.020 ;
    END
  END wbs_ack_o
  PIN wbs_adr_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 202.350 216.000 202.910 220.000 ;
    END
  END wbs_adr_i[0]
  PIN wbs_adr_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 167.390 216.000 167.950 220.000 ;
    END
  END wbs_adr_i[10]
  PIN wbs_adr_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 53.310 216.000 53.870 220.000 ;
    END
  END wbs_adr_i[11]
  PIN wbs_adr_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 130.300 4.000 131.500 ;
    END
  END wbs_adr_i[12]
  PIN wbs_adr_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 50.550 216.000 51.110 220.000 ;
    END
  END wbs_adr_i[13]
  PIN wbs_adr_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 216.000 100.380 220.000 101.580 ;
    END
  END wbs_adr_i[14]
  PIN wbs_adr_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 216.000 86.780 220.000 87.980 ;
    END
  END wbs_adr_i[15]
  PIN wbs_adr_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 106.670 0.000 107.230 4.000 ;
    END
  END wbs_adr_i[16]
  PIN wbs_adr_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 216.000 69.100 220.000 70.300 ;
    END
  END wbs_adr_i[17]
  PIN wbs_adr_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 216.000 1.100 220.000 2.300 ;
    END
  END wbs_adr_i[18]
  PIN wbs_adr_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 162.790 0.000 163.350 4.000 ;
    END
  END wbs_adr_i[19]
  PIN wbs_adr_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 192.230 216.000 192.790 220.000 ;
    END
  END wbs_adr_i[1]
  PIN wbs_adr_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 216.000 190.140 220.000 191.340 ;
    END
  END wbs_adr_i[20]
  PIN wbs_adr_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 94.710 0.000 95.270 4.000 ;
    END
  END wbs_adr_i[21]
  PIN wbs_adr_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 137.030 0.000 137.590 4.000 ;
    END
  END wbs_adr_i[22]
  PIN wbs_adr_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 206.950 0.000 207.510 4.000 ;
    END
  END wbs_adr_i[23]
  PIN wbs_adr_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 99.310 216.000 99.870 220.000 ;
    END
  END wbs_adr_i[24]
  PIN wbs_adr_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 92.870 0.000 93.430 4.000 ;
    END
  END wbs_adr_i[25]
  PIN wbs_adr_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 18.350 0.000 18.910 4.000 ;
    END
  END wbs_adr_i[26]
  PIN wbs_adr_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 137.030 216.000 137.590 220.000 ;
    END
  END wbs_adr_i[27]
  PIN wbs_adr_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 216.000 73.180 220.000 74.380 ;
    END
  END wbs_adr_i[28]
  PIN wbs_adr_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 216.000 165.660 220.000 166.860 ;
    END
  END wbs_adr_i[29]
  PIN wbs_adr_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 64.350 0.000 64.910 4.000 ;
    END
  END wbs_adr_i[2]
  PIN wbs_adr_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 211.550 216.000 212.110 220.000 ;
    END
  END wbs_adr_i[30]
  PIN wbs_adr_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 216.000 35.100 220.000 36.300 ;
    END
  END wbs_adr_i[31]
  PIN wbs_adr_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 13.340 4.000 14.540 ;
    END
  END wbs_adr_i[3]
  PIN wbs_adr_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 177.900 4.000 179.100 ;
    END
  END wbs_adr_i[4]
  PIN wbs_adr_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 127.830 0.000 128.390 4.000 ;
    END
  END wbs_adr_i[5]
  PIN wbs_adr_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 53.310 0.000 53.870 4.000 ;
    END
  END wbs_adr_i[6]
  PIN wbs_adr_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 6.540 4.000 7.740 ;
    END
  END wbs_adr_i[7]
  PIN wbs_adr_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 171.990 0.000 172.550 4.000 ;
    END
  END wbs_adr_i[8]
  PIN wbs_adr_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 217.990 0.000 218.550 4.000 ;
    END
  END wbs_adr_i[9]
  PIN wbs_cyc_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 125.070 216.000 125.630 220.000 ;
    END
  END wbs_cyc_i
  PIN wbs_dat_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 47.340 4.000 48.540 ;
    END
  END wbs_dat_i[0]
  PIN wbs_dat_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 29.390 216.000 29.950 220.000 ;
    END
  END wbs_dat_i[10]
  PIN wbs_dat_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 41.350 216.000 41.910 220.000 ;
    END
  END wbs_dat_i[11]
  PIN wbs_dat_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 33.990 216.000 34.550 220.000 ;
    END
  END wbs_dat_i[12]
  PIN wbs_dat_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 6.390 0.000 6.950 4.000 ;
    END
  END wbs_dat_i[13]
  PIN wbs_dat_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 74.540 4.000 75.740 ;
    END
  END wbs_dat_i[14]
  PIN wbs_dat_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 216.000 66.380 220.000 67.580 ;
    END
  END wbs_dat_i[15]
  PIN wbs_dat_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 99.310 0.000 99.870 4.000 ;
    END
  END wbs_dat_i[16]
  PIN wbs_dat_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 183.030 216.000 183.590 220.000 ;
    END
  END wbs_dat_i[17]
  PIN wbs_dat_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 216.000 210.540 220.000 211.740 ;
    END
  END wbs_dat_i[18]
  PIN wbs_dat_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 73.550 216.000 74.110 220.000 ;
    END
  END wbs_dat_i[19]
  PIN wbs_dat_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 150.700 4.000 151.900 ;
    END
  END wbs_dat_i[1]
  PIN wbs_dat_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 126.220 4.000 127.420 ;
    END
  END wbs_dat_i[20]
  PIN wbs_dat_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 216.000 203.740 220.000 204.940 ;
    END
  END wbs_dat_i[21]
  PIN wbs_dat_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 205.100 4.000 206.300 ;
    END
  END wbs_dat_i[22]
  PIN wbs_dat_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 216.000 138.460 220.000 139.660 ;
    END
  END wbs_dat_i[23]
  PIN wbs_dat_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 54.140 4.000 55.340 ;
    END
  END wbs_dat_i[24]
  PIN wbs_dat_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 78.620 4.000 79.820 ;
    END
  END wbs_dat_i[25]
  PIN wbs_dat_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 206.950 216.000 207.510 220.000 ;
    END
  END wbs_dat_i[26]
  PIN wbs_dat_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 102.070 216.000 102.630 220.000 ;
    END
  END wbs_dat_i[27]
  PIN wbs_dat_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 55.150 0.000 55.710 4.000 ;
    END
  END wbs_dat_i[28]
  PIN wbs_dat_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 216.000 93.580 220.000 94.780 ;
    END
  END wbs_dat_i[29]
  PIN wbs_dat_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 143.470 0.000 144.030 4.000 ;
    END
  END wbs_dat_i[2]
  PIN wbs_dat_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 216.000 14.700 220.000 15.900 ;
    END
  END wbs_dat_i[30]
  PIN wbs_dat_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 181.980 4.000 183.180 ;
    END
  END wbs_dat_i[31]
  PIN wbs_dat_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 183.030 0.000 183.590 4.000 ;
    END
  END wbs_dat_i[3]
  PIN wbs_dat_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 27.550 0.000 28.110 4.000 ;
    END
  END wbs_dat_i[4]
  PIN wbs_dat_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 88.270 0.000 88.830 4.000 ;
    END
  END wbs_dat_i[5]
  PIN wbs_dat_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 216.000 52.780 220.000 53.980 ;
    END
  END wbs_dat_i[6]
  PIN wbs_dat_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 194.990 216.000 195.550 220.000 ;
    END
  END wbs_dat_i[7]
  PIN wbs_dat_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 216.000 172.460 220.000 173.660 ;
    END
  END wbs_dat_i[8]
  PIN wbs_dat_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 187.630 0.000 188.190 4.000 ;
    END
  END wbs_dat_i[9]
  PIN wbs_dat_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 71.820 4.000 73.020 ;
    END
  END wbs_dat_o[0]
  PIN wbs_dat_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 216.000 90.860 220.000 92.060 ;
    END
  END wbs_dat_o[10]
  PIN wbs_dat_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1.790 0.000 2.350 4.000 ;
    END
  END wbs_dat_o[11]
  PIN wbs_dat_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 216.000 183.340 220.000 184.540 ;
    END
  END wbs_dat_o[12]
  PIN wbs_dat_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 185.790 216.000 186.350 220.000 ;
    END
  END wbs_dat_o[13]
  PIN wbs_dat_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 199.590 0.000 200.150 4.000 ;
    END
  END wbs_dat_o[14]
  PIN wbs_dat_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 178.430 216.000 178.990 220.000 ;
    END
  END wbs_dat_o[15]
  PIN wbs_dat_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 99.020 4.000 100.220 ;
    END
  END wbs_dat_o[16]
  PIN wbs_dat_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 108.540 4.000 109.740 ;
    END
  END wbs_dat_o[17]
  PIN wbs_dat_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 120.470 0.000 121.030 4.000 ;
    END
  END wbs_dat_o[18]
  PIN wbs_dat_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT -0.050 0.000 0.510 4.000 ;
    END
  END wbs_dat_o[19]
  PIN wbs_dat_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 141.630 0.000 142.190 4.000 ;
    END
  END wbs_dat_o[1]
  PIN wbs_dat_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 146.620 4.000 147.820 ;
    END
  END wbs_dat_o[20]
  PIN wbs_dat_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 20.140 4.000 21.340 ;
    END
  END wbs_dat_o[21]
  PIN wbs_dat_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 94.710 216.000 95.270 220.000 ;
    END
  END wbs_dat_o[22]
  PIN wbs_dat_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 105.820 4.000 107.020 ;
    END
  END wbs_dat_o[23]
  PIN wbs_dat_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 36.750 0.000 37.310 4.000 ;
    END
  END wbs_dat_o[24]
  PIN wbs_dat_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 13.750 0.000 14.310 4.000 ;
    END
  END wbs_dat_o[25]
  PIN wbs_dat_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 138.870 216.000 139.430 220.000 ;
    END
  END wbs_dat_o[26]
  PIN wbs_dat_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 97.470 216.000 98.030 220.000 ;
    END
  END wbs_dat_o[27]
  PIN wbs_dat_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 97.470 0.000 98.030 4.000 ;
    END
  END wbs_dat_o[28]
  PIN wbs_dat_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 169.230 216.000 169.790 220.000 ;
    END
  END wbs_dat_o[29]
  PIN wbs_dat_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 216.000 17.420 220.000 18.620 ;
    END
  END wbs_dat_o[2]
  PIN wbs_dat_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 188.780 4.000 189.980 ;
    END
  END wbs_dat_o[30]
  PIN wbs_dat_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 216.000 152.060 220.000 153.260 ;
    END
  END wbs_dat_o[31]
  PIN wbs_dat_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 39.510 0.000 40.070 4.000 ;
    END
  END wbs_dat_o[3]
  PIN wbs_dat_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 68.950 0.000 69.510 4.000 ;
    END
  END wbs_dat_o[4]
  PIN wbs_dat_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 108.510 0.000 109.070 4.000 ;
    END
  END wbs_dat_o[5]
  PIN wbs_dat_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 216.000 145.260 220.000 146.460 ;
    END
  END wbs_dat_o[6]
  PIN wbs_dat_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 111.270 0.000 111.830 4.000 ;
    END
  END wbs_dat_o[7]
  PIN wbs_dat_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 157.270 216.000 157.830 220.000 ;
    END
  END wbs_dat_o[8]
  PIN wbs_dat_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 155.430 216.000 155.990 220.000 ;
    END
  END wbs_dat_o[9]
  PIN wbs_sel_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 22.950 216.000 23.510 220.000 ;
    END
  END wbs_sel_i[0]
  PIN wbs_sel_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 55.150 216.000 55.710 220.000 ;
    END
  END wbs_sel_i[1]
  PIN wbs_sel_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 132.430 0.000 132.990 4.000 ;
    END
  END wbs_sel_i[2]
  PIN wbs_sel_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 60.940 4.000 62.140 ;
    END
  END wbs_sel_i[3]
  PIN wbs_stb_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3.630 216.000 4.190 220.000 ;
    END
  END wbs_stb_i
  PIN wbs_we_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 216.000 79.980 220.000 81.180 ;
    END
  END wbs_we_i
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 215.595 206.805 ;
      LAYER met1 ;
        RECT 0.070 3.780 216.590 206.960 ;
      LAYER met2 ;
        RECT 0.100 215.720 1.510 218.125 ;
        RECT 2.630 215.720 3.350 218.125 ;
        RECT 4.470 215.720 6.110 218.125 ;
        RECT 7.230 215.720 8.870 218.125 ;
        RECT 9.990 215.720 10.710 218.125 ;
        RECT 11.830 215.720 13.470 218.125 ;
        RECT 14.590 215.720 15.310 218.125 ;
        RECT 16.430 215.720 18.070 218.125 ;
        RECT 19.190 215.720 19.910 218.125 ;
        RECT 21.030 215.720 22.670 218.125 ;
        RECT 23.790 215.720 24.510 218.125 ;
        RECT 25.630 215.720 27.270 218.125 ;
        RECT 28.390 215.720 29.110 218.125 ;
        RECT 30.230 215.720 31.870 218.125 ;
        RECT 32.990 215.720 33.710 218.125 ;
        RECT 34.830 215.720 36.470 218.125 ;
        RECT 37.590 215.720 38.310 218.125 ;
        RECT 39.430 215.720 41.070 218.125 ;
        RECT 42.190 215.720 42.910 218.125 ;
        RECT 44.030 215.720 45.670 218.125 ;
        RECT 46.790 215.720 48.430 218.125 ;
        RECT 49.550 215.720 50.270 218.125 ;
        RECT 51.390 215.720 53.030 218.125 ;
        RECT 54.150 215.720 54.870 218.125 ;
        RECT 55.990 215.720 57.630 218.125 ;
        RECT 58.750 215.720 59.470 218.125 ;
        RECT 60.590 215.720 62.230 218.125 ;
        RECT 63.350 215.720 64.070 218.125 ;
        RECT 65.190 215.720 66.830 218.125 ;
        RECT 67.950 215.720 68.670 218.125 ;
        RECT 69.790 215.720 71.430 218.125 ;
        RECT 72.550 215.720 73.270 218.125 ;
        RECT 74.390 215.720 76.030 218.125 ;
        RECT 77.150 215.720 77.870 218.125 ;
        RECT 78.990 215.720 80.630 218.125 ;
        RECT 81.750 215.720 82.470 218.125 ;
        RECT 83.590 215.720 85.230 218.125 ;
        RECT 86.350 215.720 87.990 218.125 ;
        RECT 89.110 215.720 89.830 218.125 ;
        RECT 90.950 215.720 92.590 218.125 ;
        RECT 93.710 215.720 94.430 218.125 ;
        RECT 95.550 215.720 97.190 218.125 ;
        RECT 98.310 215.720 99.030 218.125 ;
        RECT 100.150 215.720 101.790 218.125 ;
        RECT 102.910 215.720 103.630 218.125 ;
        RECT 104.750 215.720 106.390 218.125 ;
        RECT 107.510 215.720 108.230 218.125 ;
        RECT 109.350 215.720 110.990 218.125 ;
        RECT 112.110 215.720 112.830 218.125 ;
        RECT 113.950 215.720 115.590 218.125 ;
        RECT 116.710 215.720 117.430 218.125 ;
        RECT 118.550 215.720 120.190 218.125 ;
        RECT 121.310 215.720 122.950 218.125 ;
        RECT 124.070 215.720 124.790 218.125 ;
        RECT 125.910 215.720 127.550 218.125 ;
        RECT 128.670 215.720 129.390 218.125 ;
        RECT 130.510 215.720 132.150 218.125 ;
        RECT 133.270 215.720 133.990 218.125 ;
        RECT 135.110 215.720 136.750 218.125 ;
        RECT 137.870 215.720 138.590 218.125 ;
        RECT 139.710 215.720 141.350 218.125 ;
        RECT 142.470 215.720 143.190 218.125 ;
        RECT 144.310 215.720 145.950 218.125 ;
        RECT 147.070 215.720 147.790 218.125 ;
        RECT 148.910 215.720 150.550 218.125 ;
        RECT 151.670 215.720 152.390 218.125 ;
        RECT 153.510 215.720 155.150 218.125 ;
        RECT 156.270 215.720 156.990 218.125 ;
        RECT 158.110 215.720 159.750 218.125 ;
        RECT 160.870 215.720 162.510 218.125 ;
        RECT 163.630 215.720 164.350 218.125 ;
        RECT 165.470 215.720 167.110 218.125 ;
        RECT 168.230 215.720 168.950 218.125 ;
        RECT 170.070 215.720 171.710 218.125 ;
        RECT 172.830 215.720 173.550 218.125 ;
        RECT 174.670 215.720 176.310 218.125 ;
        RECT 177.430 215.720 178.150 218.125 ;
        RECT 179.270 215.720 180.910 218.125 ;
        RECT 182.030 215.720 182.750 218.125 ;
        RECT 183.870 215.720 185.510 218.125 ;
        RECT 186.630 215.720 187.350 218.125 ;
        RECT 188.470 215.720 190.110 218.125 ;
        RECT 191.230 215.720 191.950 218.125 ;
        RECT 193.070 215.720 194.710 218.125 ;
        RECT 195.830 215.720 196.550 218.125 ;
        RECT 197.670 215.720 199.310 218.125 ;
        RECT 200.430 215.720 202.070 218.125 ;
        RECT 203.190 215.720 203.910 218.125 ;
        RECT 205.030 215.720 206.670 218.125 ;
        RECT 207.790 215.720 208.510 218.125 ;
        RECT 209.630 215.720 211.270 218.125 ;
        RECT 212.390 215.720 213.110 218.125 ;
        RECT 214.230 215.720 215.870 218.125 ;
        RECT 0.100 4.280 216.560 215.720 ;
        RECT 0.790 2.875 1.510 4.280 ;
        RECT 2.630 2.875 4.270 4.280 ;
        RECT 5.390 2.875 6.110 4.280 ;
        RECT 7.230 2.875 8.870 4.280 ;
        RECT 9.990 2.875 10.710 4.280 ;
        RECT 11.830 2.875 13.470 4.280 ;
        RECT 14.590 2.875 15.310 4.280 ;
        RECT 16.430 2.875 18.070 4.280 ;
        RECT 19.190 2.875 19.910 4.280 ;
        RECT 21.030 2.875 22.670 4.280 ;
        RECT 23.790 2.875 24.510 4.280 ;
        RECT 25.630 2.875 27.270 4.280 ;
        RECT 28.390 2.875 29.110 4.280 ;
        RECT 30.230 2.875 31.870 4.280 ;
        RECT 32.990 2.875 33.710 4.280 ;
        RECT 34.830 2.875 36.470 4.280 ;
        RECT 37.590 2.875 39.230 4.280 ;
        RECT 40.350 2.875 41.070 4.280 ;
        RECT 42.190 2.875 43.830 4.280 ;
        RECT 44.950 2.875 45.670 4.280 ;
        RECT 46.790 2.875 48.430 4.280 ;
        RECT 49.550 2.875 50.270 4.280 ;
        RECT 51.390 2.875 53.030 4.280 ;
        RECT 54.150 2.875 54.870 4.280 ;
        RECT 55.990 2.875 57.630 4.280 ;
        RECT 58.750 2.875 59.470 4.280 ;
        RECT 60.590 2.875 62.230 4.280 ;
        RECT 63.350 2.875 64.070 4.280 ;
        RECT 65.190 2.875 66.830 4.280 ;
        RECT 67.950 2.875 68.670 4.280 ;
        RECT 69.790 2.875 71.430 4.280 ;
        RECT 72.550 2.875 73.270 4.280 ;
        RECT 74.390 2.875 76.030 4.280 ;
        RECT 77.150 2.875 78.790 4.280 ;
        RECT 79.910 2.875 80.630 4.280 ;
        RECT 81.750 2.875 83.390 4.280 ;
        RECT 84.510 2.875 85.230 4.280 ;
        RECT 86.350 2.875 87.990 4.280 ;
        RECT 89.110 2.875 89.830 4.280 ;
        RECT 90.950 2.875 92.590 4.280 ;
        RECT 93.710 2.875 94.430 4.280 ;
        RECT 95.550 2.875 97.190 4.280 ;
        RECT 98.310 2.875 99.030 4.280 ;
        RECT 100.150 2.875 101.790 4.280 ;
        RECT 102.910 2.875 103.630 4.280 ;
        RECT 104.750 2.875 106.390 4.280 ;
        RECT 107.510 2.875 108.230 4.280 ;
        RECT 109.350 2.875 110.990 4.280 ;
        RECT 112.110 2.875 112.830 4.280 ;
        RECT 113.950 2.875 115.590 4.280 ;
        RECT 116.710 2.875 118.350 4.280 ;
        RECT 119.470 2.875 120.190 4.280 ;
        RECT 121.310 2.875 122.950 4.280 ;
        RECT 124.070 2.875 124.790 4.280 ;
        RECT 125.910 2.875 127.550 4.280 ;
        RECT 128.670 2.875 129.390 4.280 ;
        RECT 130.510 2.875 132.150 4.280 ;
        RECT 133.270 2.875 133.990 4.280 ;
        RECT 135.110 2.875 136.750 4.280 ;
        RECT 137.870 2.875 138.590 4.280 ;
        RECT 139.710 2.875 141.350 4.280 ;
        RECT 142.470 2.875 143.190 4.280 ;
        RECT 144.310 2.875 145.950 4.280 ;
        RECT 147.070 2.875 147.790 4.280 ;
        RECT 148.910 2.875 150.550 4.280 ;
        RECT 151.670 2.875 152.390 4.280 ;
        RECT 153.510 2.875 155.150 4.280 ;
        RECT 156.270 2.875 157.910 4.280 ;
        RECT 159.030 2.875 159.750 4.280 ;
        RECT 160.870 2.875 162.510 4.280 ;
        RECT 163.630 2.875 164.350 4.280 ;
        RECT 165.470 2.875 167.110 4.280 ;
        RECT 168.230 2.875 168.950 4.280 ;
        RECT 170.070 2.875 171.710 4.280 ;
        RECT 172.830 2.875 173.550 4.280 ;
        RECT 174.670 2.875 176.310 4.280 ;
        RECT 177.430 2.875 178.150 4.280 ;
        RECT 179.270 2.875 180.910 4.280 ;
        RECT 182.030 2.875 182.750 4.280 ;
        RECT 183.870 2.875 185.510 4.280 ;
        RECT 186.630 2.875 187.350 4.280 ;
        RECT 188.470 2.875 190.110 4.280 ;
        RECT 191.230 2.875 191.950 4.280 ;
        RECT 193.070 2.875 194.710 4.280 ;
        RECT 195.830 2.875 197.470 4.280 ;
        RECT 198.590 2.875 199.310 4.280 ;
        RECT 200.430 2.875 202.070 4.280 ;
        RECT 203.190 2.875 203.910 4.280 ;
        RECT 205.030 2.875 206.670 4.280 ;
        RECT 207.790 2.875 208.510 4.280 ;
        RECT 209.630 2.875 211.270 4.280 ;
        RECT 212.390 2.875 213.110 4.280 ;
        RECT 214.230 2.875 215.870 4.280 ;
      LAYER met3 ;
        RECT 4.000 217.580 215.600 218.105 ;
        RECT 4.400 216.940 215.600 217.580 ;
        RECT 4.400 216.220 216.000 216.940 ;
        RECT 4.400 215.580 215.600 216.220 ;
        RECT 4.000 214.220 215.600 215.580 ;
        RECT 4.000 213.500 216.000 214.220 ;
        RECT 4.400 212.140 216.000 213.500 ;
        RECT 4.400 211.500 215.600 212.140 ;
        RECT 4.000 210.780 215.600 211.500 ;
        RECT 4.400 210.140 215.600 210.780 ;
        RECT 4.400 209.420 216.000 210.140 ;
        RECT 4.400 208.780 215.600 209.420 ;
        RECT 4.000 207.420 215.600 208.780 ;
        RECT 4.000 206.700 216.000 207.420 ;
        RECT 4.400 205.340 216.000 206.700 ;
        RECT 4.400 204.700 215.600 205.340 ;
        RECT 4.000 203.980 215.600 204.700 ;
        RECT 4.400 203.340 215.600 203.980 ;
        RECT 4.400 202.620 216.000 203.340 ;
        RECT 4.400 201.980 215.600 202.620 ;
        RECT 4.000 200.620 215.600 201.980 ;
        RECT 4.000 199.900 216.000 200.620 ;
        RECT 4.400 198.540 216.000 199.900 ;
        RECT 4.400 197.900 215.600 198.540 ;
        RECT 4.000 197.180 215.600 197.900 ;
        RECT 4.400 196.540 215.600 197.180 ;
        RECT 4.400 195.820 216.000 196.540 ;
        RECT 4.400 195.180 215.600 195.820 ;
        RECT 4.000 193.820 215.600 195.180 ;
        RECT 4.000 193.100 216.000 193.820 ;
        RECT 4.400 191.740 216.000 193.100 ;
        RECT 4.400 191.100 215.600 191.740 ;
        RECT 4.000 190.380 215.600 191.100 ;
        RECT 4.400 189.740 215.600 190.380 ;
        RECT 4.400 188.380 216.000 189.740 ;
        RECT 4.000 187.660 216.000 188.380 ;
        RECT 4.000 186.300 215.600 187.660 ;
        RECT 4.400 185.660 215.600 186.300 ;
        RECT 4.400 184.940 216.000 185.660 ;
        RECT 4.400 184.300 215.600 184.940 ;
        RECT 4.000 183.580 215.600 184.300 ;
        RECT 4.400 182.940 215.600 183.580 ;
        RECT 4.400 181.580 216.000 182.940 ;
        RECT 4.000 180.860 216.000 181.580 ;
        RECT 4.000 179.500 215.600 180.860 ;
        RECT 4.400 178.860 215.600 179.500 ;
        RECT 4.400 178.140 216.000 178.860 ;
        RECT 4.400 177.500 215.600 178.140 ;
        RECT 4.000 176.780 215.600 177.500 ;
        RECT 4.400 176.140 215.600 176.780 ;
        RECT 4.400 174.780 216.000 176.140 ;
        RECT 4.000 174.060 216.000 174.780 ;
        RECT 4.000 172.700 215.600 174.060 ;
        RECT 4.400 172.060 215.600 172.700 ;
        RECT 4.400 171.340 216.000 172.060 ;
        RECT 4.400 170.700 215.600 171.340 ;
        RECT 4.000 169.340 215.600 170.700 ;
        RECT 4.000 168.620 216.000 169.340 ;
        RECT 4.400 167.260 216.000 168.620 ;
        RECT 4.400 166.620 215.600 167.260 ;
        RECT 4.000 165.900 215.600 166.620 ;
        RECT 4.400 165.260 215.600 165.900 ;
        RECT 4.400 164.540 216.000 165.260 ;
        RECT 4.400 163.900 215.600 164.540 ;
        RECT 4.000 162.540 215.600 163.900 ;
        RECT 4.000 161.820 216.000 162.540 ;
        RECT 4.400 160.460 216.000 161.820 ;
        RECT 4.400 159.820 215.600 160.460 ;
        RECT 4.000 159.100 215.600 159.820 ;
        RECT 4.400 158.460 215.600 159.100 ;
        RECT 4.400 157.740 216.000 158.460 ;
        RECT 4.400 157.100 215.600 157.740 ;
        RECT 4.000 155.740 215.600 157.100 ;
        RECT 4.000 155.020 216.000 155.740 ;
        RECT 4.400 153.660 216.000 155.020 ;
        RECT 4.400 153.020 215.600 153.660 ;
        RECT 4.000 152.300 215.600 153.020 ;
        RECT 4.400 151.660 215.600 152.300 ;
        RECT 4.400 150.940 216.000 151.660 ;
        RECT 4.400 150.300 215.600 150.940 ;
        RECT 4.000 148.940 215.600 150.300 ;
        RECT 4.000 148.220 216.000 148.940 ;
        RECT 4.400 146.860 216.000 148.220 ;
        RECT 4.400 146.220 215.600 146.860 ;
        RECT 4.000 145.500 215.600 146.220 ;
        RECT 4.400 144.860 215.600 145.500 ;
        RECT 4.400 144.140 216.000 144.860 ;
        RECT 4.400 143.500 215.600 144.140 ;
        RECT 4.000 142.140 215.600 143.500 ;
        RECT 4.000 141.420 216.000 142.140 ;
        RECT 4.400 140.060 216.000 141.420 ;
        RECT 4.400 139.420 215.600 140.060 ;
        RECT 4.000 138.700 215.600 139.420 ;
        RECT 4.400 138.060 215.600 138.700 ;
        RECT 4.400 137.340 216.000 138.060 ;
        RECT 4.400 136.700 215.600 137.340 ;
        RECT 4.000 135.340 215.600 136.700 ;
        RECT 4.000 134.620 216.000 135.340 ;
        RECT 4.400 133.260 216.000 134.620 ;
        RECT 4.400 132.620 215.600 133.260 ;
        RECT 4.000 131.900 215.600 132.620 ;
        RECT 4.400 131.260 215.600 131.900 ;
        RECT 4.400 129.900 216.000 131.260 ;
        RECT 4.000 129.180 216.000 129.900 ;
        RECT 4.000 127.820 215.600 129.180 ;
        RECT 4.400 127.180 215.600 127.820 ;
        RECT 4.400 126.460 216.000 127.180 ;
        RECT 4.400 125.820 215.600 126.460 ;
        RECT 4.000 125.100 215.600 125.820 ;
        RECT 4.400 124.460 215.600 125.100 ;
        RECT 4.400 123.100 216.000 124.460 ;
        RECT 4.000 122.380 216.000 123.100 ;
        RECT 4.000 121.020 215.600 122.380 ;
        RECT 4.400 120.380 215.600 121.020 ;
        RECT 4.400 119.660 216.000 120.380 ;
        RECT 4.400 119.020 215.600 119.660 ;
        RECT 4.000 118.300 215.600 119.020 ;
        RECT 4.400 117.660 215.600 118.300 ;
        RECT 4.400 116.300 216.000 117.660 ;
        RECT 4.000 115.580 216.000 116.300 ;
        RECT 4.000 114.220 215.600 115.580 ;
        RECT 4.400 113.580 215.600 114.220 ;
        RECT 4.400 112.860 216.000 113.580 ;
        RECT 4.400 112.220 215.600 112.860 ;
        RECT 4.000 110.860 215.600 112.220 ;
        RECT 4.000 110.140 216.000 110.860 ;
        RECT 4.400 108.780 216.000 110.140 ;
        RECT 4.400 108.140 215.600 108.780 ;
        RECT 4.000 107.420 215.600 108.140 ;
        RECT 4.400 106.780 215.600 107.420 ;
        RECT 4.400 106.060 216.000 106.780 ;
        RECT 4.400 105.420 215.600 106.060 ;
        RECT 4.000 104.060 215.600 105.420 ;
        RECT 4.000 103.340 216.000 104.060 ;
        RECT 4.400 101.980 216.000 103.340 ;
        RECT 4.400 101.340 215.600 101.980 ;
        RECT 4.000 100.620 215.600 101.340 ;
        RECT 4.400 99.980 215.600 100.620 ;
        RECT 4.400 99.260 216.000 99.980 ;
        RECT 4.400 98.620 215.600 99.260 ;
        RECT 4.000 97.260 215.600 98.620 ;
        RECT 4.000 96.540 216.000 97.260 ;
        RECT 4.400 95.180 216.000 96.540 ;
        RECT 4.400 94.540 215.600 95.180 ;
        RECT 4.000 93.820 215.600 94.540 ;
        RECT 4.400 93.180 215.600 93.820 ;
        RECT 4.400 92.460 216.000 93.180 ;
        RECT 4.400 91.820 215.600 92.460 ;
        RECT 4.000 90.460 215.600 91.820 ;
        RECT 4.000 89.740 216.000 90.460 ;
        RECT 4.400 88.380 216.000 89.740 ;
        RECT 4.400 87.740 215.600 88.380 ;
        RECT 4.000 87.020 215.600 87.740 ;
        RECT 4.400 86.380 215.600 87.020 ;
        RECT 4.400 85.660 216.000 86.380 ;
        RECT 4.400 85.020 215.600 85.660 ;
        RECT 4.000 83.660 215.600 85.020 ;
        RECT 4.000 82.940 216.000 83.660 ;
        RECT 4.400 81.580 216.000 82.940 ;
        RECT 4.400 80.940 215.600 81.580 ;
        RECT 4.000 80.220 215.600 80.940 ;
        RECT 4.400 79.580 215.600 80.220 ;
        RECT 4.400 78.860 216.000 79.580 ;
        RECT 4.400 78.220 215.600 78.860 ;
        RECT 4.000 76.860 215.600 78.220 ;
        RECT 4.000 76.140 216.000 76.860 ;
        RECT 4.400 74.780 216.000 76.140 ;
        RECT 4.400 74.140 215.600 74.780 ;
        RECT 4.000 73.420 215.600 74.140 ;
        RECT 4.400 72.780 215.600 73.420 ;
        RECT 4.400 71.420 216.000 72.780 ;
        RECT 4.000 70.700 216.000 71.420 ;
        RECT 4.000 69.340 215.600 70.700 ;
        RECT 4.400 68.700 215.600 69.340 ;
        RECT 4.400 67.980 216.000 68.700 ;
        RECT 4.400 67.340 215.600 67.980 ;
        RECT 4.000 66.620 215.600 67.340 ;
        RECT 4.400 65.980 215.600 66.620 ;
        RECT 4.400 64.620 216.000 65.980 ;
        RECT 4.000 63.900 216.000 64.620 ;
        RECT 4.000 62.540 215.600 63.900 ;
        RECT 4.400 61.900 215.600 62.540 ;
        RECT 4.400 61.180 216.000 61.900 ;
        RECT 4.400 60.540 215.600 61.180 ;
        RECT 4.000 59.820 215.600 60.540 ;
        RECT 4.400 59.180 215.600 59.820 ;
        RECT 4.400 57.820 216.000 59.180 ;
        RECT 4.000 57.100 216.000 57.820 ;
        RECT 4.000 55.740 215.600 57.100 ;
        RECT 4.400 55.100 215.600 55.740 ;
        RECT 4.400 54.380 216.000 55.100 ;
        RECT 4.400 53.740 215.600 54.380 ;
        RECT 4.000 52.380 215.600 53.740 ;
        RECT 4.000 51.660 216.000 52.380 ;
        RECT 4.400 50.300 216.000 51.660 ;
        RECT 4.400 49.660 215.600 50.300 ;
        RECT 4.000 48.940 215.600 49.660 ;
        RECT 4.400 48.300 215.600 48.940 ;
        RECT 4.400 47.580 216.000 48.300 ;
        RECT 4.400 46.940 215.600 47.580 ;
        RECT 4.000 45.580 215.600 46.940 ;
        RECT 4.000 44.860 216.000 45.580 ;
        RECT 4.400 43.500 216.000 44.860 ;
        RECT 4.400 42.860 215.600 43.500 ;
        RECT 4.000 42.140 215.600 42.860 ;
        RECT 4.400 41.500 215.600 42.140 ;
        RECT 4.400 40.780 216.000 41.500 ;
        RECT 4.400 40.140 215.600 40.780 ;
        RECT 4.000 38.780 215.600 40.140 ;
        RECT 4.000 38.060 216.000 38.780 ;
        RECT 4.400 36.700 216.000 38.060 ;
        RECT 4.400 36.060 215.600 36.700 ;
        RECT 4.000 35.340 215.600 36.060 ;
        RECT 4.400 34.700 215.600 35.340 ;
        RECT 4.400 33.980 216.000 34.700 ;
        RECT 4.400 33.340 215.600 33.980 ;
        RECT 4.000 31.980 215.600 33.340 ;
        RECT 4.000 31.260 216.000 31.980 ;
        RECT 4.400 29.900 216.000 31.260 ;
        RECT 4.400 29.260 215.600 29.900 ;
        RECT 4.000 28.540 215.600 29.260 ;
        RECT 4.400 27.900 215.600 28.540 ;
        RECT 4.400 27.180 216.000 27.900 ;
        RECT 4.400 26.540 215.600 27.180 ;
        RECT 4.000 25.180 215.600 26.540 ;
        RECT 4.000 24.460 216.000 25.180 ;
        RECT 4.400 23.100 216.000 24.460 ;
        RECT 4.400 22.460 215.600 23.100 ;
        RECT 4.000 21.740 215.600 22.460 ;
        RECT 4.400 21.100 215.600 21.740 ;
        RECT 4.400 19.740 216.000 21.100 ;
        RECT 4.000 19.020 216.000 19.740 ;
        RECT 4.000 17.660 215.600 19.020 ;
        RECT 4.400 17.020 215.600 17.660 ;
        RECT 4.400 16.300 216.000 17.020 ;
        RECT 4.400 15.660 215.600 16.300 ;
        RECT 4.000 14.940 215.600 15.660 ;
        RECT 4.400 14.300 215.600 14.940 ;
        RECT 4.400 12.940 216.000 14.300 ;
        RECT 4.000 12.220 216.000 12.940 ;
        RECT 4.000 10.860 215.600 12.220 ;
        RECT 4.400 10.220 215.600 10.860 ;
        RECT 4.400 9.500 216.000 10.220 ;
        RECT 4.400 8.860 215.600 9.500 ;
        RECT 4.000 8.140 215.600 8.860 ;
        RECT 4.400 7.500 215.600 8.140 ;
        RECT 4.400 6.140 216.000 7.500 ;
        RECT 4.000 5.420 216.000 6.140 ;
        RECT 4.000 4.060 215.600 5.420 ;
        RECT 4.400 3.420 215.600 4.060 ;
        RECT 4.400 2.895 216.000 3.420 ;
  END
END wrapped_asic_watch
END LIBRARY

