VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO wrapped_asic_watch
  CLASS BLOCK ;
  FOREIGN wrapped_asic_watch ;
  ORIGIN 0.000 0.000 ;
  SIZE 300.000 BY 300.000 ;
  PIN active
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 24.790 296.000 25.350 300.000 ;
    END
  END active
  PIN io_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 79.990 0.000 80.550 4.000 ;
    END
  END io_in[0]
  PIN io_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 185.790 296.000 186.350 300.000 ;
    END
  END io_in[10]
  PIN io_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 43.190 296.000 43.750 300.000 ;
    END
  END io_in[11]
  PIN io_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 241.820 300.000 243.020 ;
    END
  END io_in[12]
  PIN io_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 122.310 0.000 122.870 4.000 ;
    END
  END io_in[13]
  PIN io_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 137.950 296.000 138.510 300.000 ;
    END
  END io_in[14]
  PIN io_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 256.780 300.000 257.980 ;
    END
  END io_in[15]
  PIN io_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 278.710 0.000 279.270 4.000 ;
    END
  END io_in[16]
  PIN io_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 95.630 296.000 96.190 300.000 ;
    END
  END io_in[17]
  PIN io_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 104.830 296.000 105.390 300.000 ;
    END
  END io_in[18]
  PIN io_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 222.590 0.000 223.150 4.000 ;
    END
  END io_in[19]
  PIN io_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 118.060 4.000 119.260 ;
    END
  END io_in[1]
  PIN io_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 209.180 4.000 210.380 ;
    END
  END io_in[20]
  PIN io_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 139.820 4.000 141.020 ;
    END
  END io_in[21]
  PIN io_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 52.780 300.000 53.980 ;
    END
  END io_in[22]
  PIN io_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 91.030 296.000 91.590 300.000 ;
    END
  END io_in[23]
  PIN io_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 76.310 296.000 76.870 300.000 ;
    END
  END io_in[24]
  PIN io_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 194.070 0.000 194.630 4.000 ;
    END
  END io_in[25]
  PIN io_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 189.470 0.000 190.030 4.000 ;
    END
  END io_in[26]
  PIN io_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 17.420 300.000 18.620 ;
    END
  END io_in[27]
  PIN io_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 170.150 0.000 170.710 4.000 ;
    END
  END io_in[28]
  PIN io_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 298.950 296.000 299.510 300.000 ;
    END
  END io_in[29]
  PIN io_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 84.590 0.000 85.150 4.000 ;
    END
  END io_in[2]
  PIN io_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 81.340 300.000 82.540 ;
    END
  END io_in[30]
  PIN io_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 14.670 296.000 15.230 300.000 ;
    END
  END io_in[31]
  PIN io_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 160.950 0.000 161.510 4.000 ;
    END
  END io_in[32]
  PIN io_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 188.780 4.000 189.980 ;
    END
  END io_in[33]
  PIN io_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 238.230 296.000 238.790 300.000 ;
    END
  END io_in[34]
  PIN io_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 265.830 296.000 266.390 300.000 ;
    END
  END io_in[35]
  PIN io_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 165.660 300.000 166.860 ;
    END
  END io_in[36]
  PIN io_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 271.350 296.000 271.910 300.000 ;
    END
  END io_in[37]
  PIN io_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 190.390 296.000 190.950 300.000 ;
    END
  END io_in[3]
  PIN io_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 157.500 300.000 158.700 ;
    END
  END io_in[4]
  PIN io_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 283.980 300.000 285.180 ;
    END
  END io_in[5]
  PIN io_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 222.780 4.000 223.980 ;
    END
  END io_in[6]
  PIN io_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 153.420 4.000 154.620 ;
    END
  END io_in[7]
  PIN io_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 179.260 300.000 180.460 ;
    END
  END io_in[8]
  PIN io_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 86.430 296.000 86.990 300.000 ;
    END
  END io_in[9]
  PIN io_oeb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 137.030 0.000 137.590 4.000 ;
    END
  END io_oeb[0]
  PIN io_oeb[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 124.860 4.000 126.060 ;
    END
  END io_oeb[10]
  PIN io_oeb[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 143.900 300.000 145.100 ;
    END
  END io_oeb[11]
  PIN io_oeb[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 45.980 300.000 47.180 ;
    END
  END io_oeb[12]
  PIN io_oeb[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 39.180 300.000 40.380 ;
    END
  END io_oeb[13]
  PIN io_oeb[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 33.740 4.000 34.940 ;
    END
  END io_oeb[14]
  PIN io_oeb[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 114.950 296.000 115.510 300.000 ;
    END
  END io_oeb[15]
  PIN io_oeb[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 269.510 0.000 270.070 4.000 ;
    END
  END io_oeb[16]
  PIN io_oeb[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 70.790 0.000 71.350 4.000 ;
    END
  END io_oeb[17]
  PIN io_oeb[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 228.110 296.000 228.670 300.000 ;
    END
  END io_oeb[18]
  PIN io_oeb[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 119.550 296.000 120.110 300.000 ;
    END
  END io_oeb[19]
  PIN io_oeb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 203.270 0.000 203.830 4.000 ;
    END
  END io_oeb[1]
  PIN io_oeb[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 94.940 300.000 96.140 ;
    END
  END io_oeb[20]
  PIN io_oeb[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 53.310 296.000 53.870 300.000 ;
    END
  END io_oeb[21]
  PIN io_oeb[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 27.550 0.000 28.110 4.000 ;
    END
  END io_oeb[22]
  PIN io_oeb[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 171.070 296.000 171.630 300.000 ;
    END
  END io_oeb[23]
  PIN io_oeb[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 176.590 296.000 177.150 300.000 ;
    END
  END io_oeb[24]
  PIN io_oeb[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 245.590 0.000 246.150 4.000 ;
    END
  END io_oeb[25]
  PIN io_oeb[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 221.420 300.000 222.620 ;
    END
  END io_oeb[26]
  PIN io_oeb[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 194.990 296.000 195.550 300.000 ;
    END
  END io_oeb[27]
  PIN io_oeb[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 217.070 0.000 217.630 4.000 ;
    END
  END io_oeb[28]
  PIN io_oeb[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 172.460 300.000 173.660 ;
    END
  END io_oeb[29]
  PIN io_oeb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 256.630 296.000 257.190 300.000 ;
    END
  END io_oeb[2]
  PIN io_oeb[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 57.910 296.000 58.470 300.000 ;
    END
  END io_oeb[30]
  PIN io_oeb[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 212.470 0.000 213.030 4.000 ;
    END
  END io_oeb[31]
  PIN io_oeb[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 180.620 4.000 181.820 ;
    END
  END io_oeb[32]
  PIN io_oeb[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 251.110 0.000 251.670 4.000 ;
    END
  END io_oeb[33]
  PIN io_oeb[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 100.230 296.000 100.790 300.000 ;
    END
  END io_oeb[34]
  PIN io_oeb[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 160.220 4.000 161.420 ;
    END
  END io_oeb[35]
  PIN io_oeb[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 82.700 4.000 83.900 ;
    END
  END io_oeb[36]
  PIN io_oeb[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 131.660 4.000 132.860 ;
    END
  END io_oeb[37]
  PIN io_oeb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 132.430 0.000 132.990 4.000 ;
    END
  END io_oeb[3]
  PIN io_oeb[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 260.310 0.000 260.870 4.000 ;
    END
  END io_oeb[4]
  PIN io_oeb[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 237.740 4.000 238.940 ;
    END
  END io_oeb[5]
  PIN io_oeb[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 67.740 300.000 68.940 ;
    END
  END io_oeb[6]
  PIN io_oeb[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 109.430 296.000 109.990 300.000 ;
    END
  END io_oeb[7]
  PIN io_oeb[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 22.950 0.000 23.510 4.000 ;
    END
  END io_oeb[8]
  PIN io_oeb[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 56.070 0.000 56.630 4.000 ;
    END
  END io_oeb[9]
  PIN io_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 277.180 300.000 278.380 ;
    END
  END io_out[0]
  PIN io_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 137.100 300.000 138.300 ;
    END
  END io_out[10]
  PIN io_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 20.140 4.000 21.340 ;
    END
  END io_out[11]
  PIN io_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 55.500 4.000 56.700 ;
    END
  END io_out[12]
  PIN io_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 207.870 0.000 208.430 4.000 ;
    END
  END io_out[13]
  PIN io_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 228.220 300.000 229.420 ;
    END
  END io_out[14]
  PIN io_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.870 296.000 1.430 300.000 ;
    END
  END io_out[15]
  PIN io_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 130.300 300.000 131.500 ;
    END
  END io_out[16]
  PIN io_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 280.550 296.000 281.110 300.000 ;
    END
  END io_out[17]
  PIN io_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 240.990 0.000 241.550 4.000 ;
    END
  END io_out[18]
  PIN io_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 173.820 4.000 175.020 ;
    END
  END io_out[19]
  PIN io_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 214.310 296.000 214.870 300.000 ;
    END
  END io_out[1]
  PIN io_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 252.030 296.000 252.590 300.000 ;
    END
  END io_out[20]
  PIN io_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 293.500 4.000 294.700 ;
    END
  END io_out[21]
  PIN io_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 165.550 0.000 166.110 4.000 ;
    END
  END io_out[22]
  PIN io_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 101.740 300.000 102.940 ;
    END
  END io_out[23]
  PIN io_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 141.630 0.000 142.190 4.000 ;
    END
  END io_out[24]
  PIN io_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 232.710 296.000 233.270 300.000 ;
    END
  END io_out[25]
  PIN io_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 40.540 4.000 41.740 ;
    END
  END io_out[26]
  PIN io_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 242.830 296.000 243.390 300.000 ;
    END
  END io_out[27]
  PIN io_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 89.190 0.000 89.750 4.000 ;
    END
  END io_out[28]
  PIN io_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 264.910 0.000 265.470 4.000 ;
    END
  END io_out[29]
  PIN io_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 37.670 0.000 38.230 4.000 ;
    END
  END io_out[2]
  PIN io_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 48.700 4.000 49.900 ;
    END
  END io_out[30]
  PIN io_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 104.460 4.000 105.660 ;
    END
  END io_out[31]
  PIN io_out[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 29.390 296.000 29.950 300.000 ;
    END
  END io_out[32]
  PIN io_out[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 293.430 0.000 293.990 4.000 ;
    END
  END io_out[33]
  PIN io_out[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 235.020 300.000 236.220 ;
    END
  END io_out[34]
  PIN io_out[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 214.620 300.000 215.820 ;
    END
  END io_out[35]
  PIN io_out[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 124.150 296.000 124.710 300.000 ;
    END
  END io_out[36]
  PIN io_out[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 263.580 300.000 264.780 ;
    END
  END io_out[37]
  PIN io_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 10.070 296.000 10.630 300.000 ;
    END
  END io_out[3]
  PIN io_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 150.700 300.000 151.900 ;
    END
  END io_out[4]
  PIN io_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 161.870 296.000 162.430 300.000 ;
    END
  END io_out[5]
  PIN io_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 289.750 296.000 290.310 300.000 ;
    END
  END io_out[6]
  PIN io_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 146.620 4.000 147.820 ;
    END
  END io_out[7]
  PIN io_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 99.310 0.000 99.870 4.000 ;
    END
  END io_out[8]
  PIN io_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 111.260 4.000 112.460 ;
    END
  END io_out[9]
  PIN la1_data_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 298.030 0.000 298.590 4.000 ;
    END
  END la1_data_in[0]
  PIN la1_data_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 113.110 0.000 113.670 4.000 ;
    END
  END la1_data_in[10]
  PIN la1_data_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 288.830 0.000 289.390 4.000 ;
    END
  END la1_data_in[11]
  PIN la1_data_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 271.740 4.000 272.940 ;
    END
  END la1_data_in[12]
  PIN la1_data_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 174.750 0.000 175.310 4.000 ;
    END
  END la1_data_in[13]
  PIN la1_data_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 97.660 4.000 98.860 ;
    END
  END la1_data_in[14]
  PIN la1_data_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 128.750 296.000 129.310 300.000 ;
    END
  END la1_data_in[15]
  PIN la1_data_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 204.190 296.000 204.750 300.000 ;
    END
  END la1_data_in[16]
  PIN la1_data_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 166.470 296.000 167.030 300.000 ;
    END
  END la1_data_in[17]
  PIN la1_data_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 227.190 0.000 227.750 4.000 ;
    END
  END la1_data_in[18]
  PIN la1_data_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 133.350 296.000 133.910 300.000 ;
    END
  END la1_data_in[19]
  PIN la1_data_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 103.910 0.000 104.470 4.000 ;
    END
  END la1_data_in[1]
  PIN la1_data_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 264.940 4.000 266.140 ;
    END
  END la1_data_in[20]
  PIN la1_data_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 294.350 296.000 294.910 300.000 ;
    END
  END la1_data_in[21]
  PIN la1_data_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 3.820 300.000 5.020 ;
    END
  END la1_data_in[22]
  PIN la1_data_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 6.540 4.000 7.740 ;
    END
  END la1_data_in[23]
  PIN la1_data_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 75.390 0.000 75.950 4.000 ;
    END
  END la1_data_in[24]
  PIN la1_data_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 279.900 4.000 281.100 ;
    END
  END la1_data_in[25]
  PIN la1_data_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 274.110 0.000 274.670 4.000 ;
    END
  END la1_data_in[26]
  PIN la1_data_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 150.830 0.000 151.390 4.000 ;
    END
  END la1_data_in[27]
  PIN la1_data_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 244.540 4.000 245.740 ;
    END
  END la1_data_in[28]
  PIN la1_data_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 47.790 296.000 48.350 300.000 ;
    END
  END la1_data_in[29]
  PIN la1_data_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 60.670 0.000 61.230 4.000 ;
    END
  END la1_data_in[2]
  PIN la1_data_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 9.150 0.000 9.710 4.000 ;
    END
  END la1_data_in[30]
  PIN la1_data_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 198.670 0.000 199.230 4.000 ;
    END
  END la1_data_in[31]
  PIN la1_data_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 229.580 4.000 230.780 ;
    END
  END la1_data_in[3]
  PIN la1_data_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 261.230 296.000 261.790 300.000 ;
    END
  END la1_data_in[4]
  PIN la1_data_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 116.700 300.000 117.900 ;
    END
  END la1_data_in[5]
  PIN la1_data_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 143.470 296.000 144.030 300.000 ;
    END
  END la1_data_in[6]
  PIN la1_data_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 167.020 4.000 168.220 ;
    END
  END la1_data_in[7]
  PIN la1_data_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 148.070 296.000 148.630 300.000 ;
    END
  END la1_data_in[8]
  PIN la1_data_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 251.340 4.000 252.540 ;
    END
  END la1_data_in[9]
  PIN la1_data_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 42.270 0.000 42.830 4.000 ;
    END
  END la1_data_out[0]
  PIN la1_data_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 25.580 300.000 26.780 ;
    END
  END la1_data_out[10]
  PIN la1_data_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 117.710 0.000 118.270 4.000 ;
    END
  END la1_data_out[11]
  PIN la1_data_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 270.380 300.000 271.580 ;
    END
  END la1_data_out[12]
  PIN la1_data_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 67.110 296.000 67.670 300.000 ;
    END
  END la1_data_out[13]
  PIN la1_data_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 181.190 296.000 181.750 300.000 ;
    END
  END la1_data_out[14]
  PIN la1_data_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 13.340 4.000 14.540 ;
    END
  END la1_data_out[15]
  PIN la1_data_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 59.580 300.000 60.780 ;
    END
  END la1_data_out[16]
  PIN la1_data_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 199.660 300.000 200.860 ;
    END
  END la1_data_out[17]
  PIN la1_data_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 71.710 296.000 72.270 300.000 ;
    END
  END la1_data_out[18]
  PIN la1_data_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 123.500 300.000 124.700 ;
    END
  END la1_data_out[19]
  PIN la1_data_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 20.190 296.000 20.750 300.000 ;
    END
  END la1_data_out[1]
  PIN la1_data_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 75.900 4.000 77.100 ;
    END
  END la1_data_out[20]
  PIN la1_data_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 248.620 300.000 249.820 ;
    END
  END la1_data_out[21]
  PIN la1_data_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 199.590 296.000 200.150 300.000 ;
    END
  END la1_data_out[22]
  PIN la1_data_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 66.190 0.000 66.750 4.000 ;
    END
  END la1_data_out[23]
  PIN la1_data_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 74.540 300.000 75.740 ;
    END
  END la1_data_out[24]
  PIN la1_data_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 26.940 4.000 28.140 ;
    END
  END la1_data_out[25]
  PIN la1_data_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 284.230 0.000 284.790 4.000 ;
    END
  END la1_data_out[26]
  PIN la1_data_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 33.990 296.000 34.550 300.000 ;
    END
  END la1_data_out[27]
  PIN la1_data_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 231.790 0.000 232.350 4.000 ;
    END
  END la1_data_out[28]
  PIN la1_data_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 33.070 0.000 33.630 4.000 ;
    END
  END la1_data_out[29]
  PIN la1_data_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 108.510 0.000 109.070 4.000 ;
    END
  END la1_data_out[2]
  PIN la1_data_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 32.380 300.000 33.580 ;
    END
  END la1_data_out[30]
  PIN la1_data_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 290.780 300.000 291.980 ;
    END
  END la1_data_out[31]
  PIN la1_data_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 69.100 4.000 70.300 ;
    END
  END la1_data_out[3]
  PIN la1_data_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 236.390 0.000 236.950 4.000 ;
    END
  END la1_data_out[4]
  PIN la1_data_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 18.350 0.000 18.910 4.000 ;
    END
  END la1_data_out[5]
  PIN la1_data_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 88.140 300.000 89.340 ;
    END
  END la1_data_out[6]
  PIN la1_data_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 4.550 0.000 5.110 4.000 ;
    END
  END la1_data_out[7]
  PIN la1_data_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 207.820 300.000 209.020 ;
    END
  END la1_data_out[8]
  PIN la1_data_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 285.150 296.000 285.710 300.000 ;
    END
  END la1_data_out[9]
  PIN la1_oenb[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 255.710 0.000 256.270 4.000 ;
    END
  END la1_oenb[0]
  PIN la1_oenb[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 275.950 296.000 276.510 300.000 ;
    END
  END la1_oenb[10]
  PIN la1_oenb[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 202.380 4.000 203.580 ;
    END
  END la1_oenb[11]
  PIN la1_oenb[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 215.980 4.000 217.180 ;
    END
  END la1_oenb[12]
  PIN la1_oenb[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 155.430 0.000 155.990 4.000 ;
    END
  END la1_oenb[13]
  PIN la1_oenb[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT -0.050 0.000 0.510 4.000 ;
    END
  END la1_oenb[14]
  PIN la1_oenb[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 183.950 0.000 184.510 4.000 ;
    END
  END la1_oenb[15]
  PIN la1_oenb[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 258.140 4.000 259.340 ;
    END
  END la1_oenb[16]
  PIN la1_oenb[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 62.510 296.000 63.070 300.000 ;
    END
  END la1_oenb[17]
  PIN la1_oenb[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 157.270 296.000 157.830 300.000 ;
    END
  END la1_oenb[18]
  PIN la1_oenb[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 195.580 4.000 196.780 ;
    END
  END la1_oenb[19]
  PIN la1_oenb[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 46.870 0.000 47.430 4.000 ;
    END
  END la1_oenb[1]
  PIN la1_oenb[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 13.750 0.000 14.310 4.000 ;
    END
  END la1_oenb[20]
  PIN la1_oenb[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 209.710 296.000 210.270 300.000 ;
    END
  END la1_oenb[21]
  PIN la1_oenb[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 152.670 296.000 153.230 300.000 ;
    END
  END la1_oenb[22]
  PIN la1_oenb[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 127.830 0.000 128.390 4.000 ;
    END
  END la1_oenb[23]
  PIN la1_oenb[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 247.430 296.000 247.990 300.000 ;
    END
  END la1_oenb[24]
  PIN la1_oenb[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 10.620 300.000 11.820 ;
    END
  END la1_oenb[25]
  PIN la1_oenb[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 286.700 4.000 287.900 ;
    END
  END la1_oenb[26]
  PIN la1_oenb[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 192.860 300.000 194.060 ;
    END
  END la1_oenb[27]
  PIN la1_oenb[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 51.470 0.000 52.030 4.000 ;
    END
  END la1_oenb[28]
  PIN la1_oenb[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 94.710 0.000 95.270 4.000 ;
    END
  END la1_oenb[29]
  PIN la1_oenb[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 62.300 4.000 63.500 ;
    END
  END la1_oenb[2]
  PIN la1_oenb[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 186.060 300.000 187.260 ;
    END
  END la1_oenb[30]
  PIN la1_oenb[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 146.230 0.000 146.790 4.000 ;
    END
  END la1_oenb[31]
  PIN la1_oenb[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 223.510 296.000 224.070 300.000 ;
    END
  END la1_oenb[3]
  PIN la1_oenb[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 218.910 296.000 219.470 300.000 ;
    END
  END la1_oenb[4]
  PIN la1_oenb[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 38.590 296.000 39.150 300.000 ;
    END
  END la1_oenb[5]
  PIN la1_oenb[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 81.830 296.000 82.390 300.000 ;
    END
  END la1_oenb[6]
  PIN la1_oenb[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 179.350 0.000 179.910 4.000 ;
    END
  END la1_oenb[7]
  PIN la1_oenb[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 89.500 4.000 90.700 ;
    END
  END la1_oenb[8]
  PIN la1_oenb[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 5.470 296.000 6.030 300.000 ;
    END
  END la1_oenb[9]
  PIN vccd1
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 288.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 288.560 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 288.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 288.560 ;
    END
  END vssd1
  PIN wb_clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 108.540 300.000 109.740 ;
    END
  END wb_clk_i
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 296.095 288.405 ;
      LAYER met1 ;
        RECT 0.990 10.640 296.155 288.560 ;
      LAYER met2 ;
        RECT 1.710 295.720 5.190 296.210 ;
        RECT 6.310 295.720 9.790 296.210 ;
        RECT 10.910 295.720 14.390 296.210 ;
        RECT 15.510 295.720 19.910 296.210 ;
        RECT 21.030 295.720 24.510 296.210 ;
        RECT 25.630 295.720 29.110 296.210 ;
        RECT 30.230 295.720 33.710 296.210 ;
        RECT 34.830 295.720 38.310 296.210 ;
        RECT 39.430 295.720 42.910 296.210 ;
        RECT 44.030 295.720 47.510 296.210 ;
        RECT 48.630 295.720 53.030 296.210 ;
        RECT 54.150 295.720 57.630 296.210 ;
        RECT 58.750 295.720 62.230 296.210 ;
        RECT 63.350 295.720 66.830 296.210 ;
        RECT 67.950 295.720 71.430 296.210 ;
        RECT 72.550 295.720 76.030 296.210 ;
        RECT 77.150 295.720 81.550 296.210 ;
        RECT 82.670 295.720 86.150 296.210 ;
        RECT 87.270 295.720 90.750 296.210 ;
        RECT 91.870 295.720 95.350 296.210 ;
        RECT 96.470 295.720 99.950 296.210 ;
        RECT 101.070 295.720 104.550 296.210 ;
        RECT 105.670 295.720 109.150 296.210 ;
        RECT 110.270 295.720 114.670 296.210 ;
        RECT 115.790 295.720 119.270 296.210 ;
        RECT 120.390 295.720 123.870 296.210 ;
        RECT 124.990 295.720 128.470 296.210 ;
        RECT 129.590 295.720 133.070 296.210 ;
        RECT 134.190 295.720 137.670 296.210 ;
        RECT 138.790 295.720 143.190 296.210 ;
        RECT 144.310 295.720 147.790 296.210 ;
        RECT 148.910 295.720 152.390 296.210 ;
        RECT 153.510 295.720 156.990 296.210 ;
        RECT 158.110 295.720 161.590 296.210 ;
        RECT 162.710 295.720 166.190 296.210 ;
        RECT 167.310 295.720 170.790 296.210 ;
        RECT 171.910 295.720 176.310 296.210 ;
        RECT 177.430 295.720 180.910 296.210 ;
        RECT 182.030 295.720 185.510 296.210 ;
        RECT 186.630 295.720 190.110 296.210 ;
        RECT 191.230 295.720 194.710 296.210 ;
        RECT 195.830 295.720 199.310 296.210 ;
        RECT 200.430 295.720 203.910 296.210 ;
        RECT 205.030 295.720 209.430 296.210 ;
        RECT 210.550 295.720 214.030 296.210 ;
        RECT 215.150 295.720 218.630 296.210 ;
        RECT 219.750 295.720 223.230 296.210 ;
        RECT 224.350 295.720 227.830 296.210 ;
        RECT 228.950 295.720 232.430 296.210 ;
        RECT 233.550 295.720 237.950 296.210 ;
        RECT 239.070 295.720 242.550 296.210 ;
        RECT 243.670 295.720 247.150 296.210 ;
        RECT 248.270 295.720 251.750 296.210 ;
        RECT 252.870 295.720 256.350 296.210 ;
        RECT 257.470 295.720 260.950 296.210 ;
        RECT 262.070 295.720 265.550 296.210 ;
        RECT 266.670 295.720 271.070 296.210 ;
        RECT 272.190 295.720 275.670 296.210 ;
        RECT 276.790 295.720 280.270 296.210 ;
        RECT 281.390 295.720 284.870 296.210 ;
        RECT 285.990 295.720 289.470 296.210 ;
        RECT 290.590 295.720 293.840 296.210 ;
        RECT 1.020 4.280 293.840 295.720 ;
        RECT 1.020 4.000 4.270 4.280 ;
        RECT 5.390 4.000 8.870 4.280 ;
        RECT 9.990 4.000 13.470 4.280 ;
        RECT 14.590 4.000 18.070 4.280 ;
        RECT 19.190 4.000 22.670 4.280 ;
        RECT 23.790 4.000 27.270 4.280 ;
        RECT 28.390 4.000 32.790 4.280 ;
        RECT 33.910 4.000 37.390 4.280 ;
        RECT 38.510 4.000 41.990 4.280 ;
        RECT 43.110 4.000 46.590 4.280 ;
        RECT 47.710 4.000 51.190 4.280 ;
        RECT 52.310 4.000 55.790 4.280 ;
        RECT 56.910 4.000 60.390 4.280 ;
        RECT 61.510 4.000 65.910 4.280 ;
        RECT 67.030 4.000 70.510 4.280 ;
        RECT 71.630 4.000 75.110 4.280 ;
        RECT 76.230 4.000 79.710 4.280 ;
        RECT 80.830 4.000 84.310 4.280 ;
        RECT 85.430 4.000 88.910 4.280 ;
        RECT 90.030 4.000 94.430 4.280 ;
        RECT 95.550 4.000 99.030 4.280 ;
        RECT 100.150 4.000 103.630 4.280 ;
        RECT 104.750 4.000 108.230 4.280 ;
        RECT 109.350 4.000 112.830 4.280 ;
        RECT 113.950 4.000 117.430 4.280 ;
        RECT 118.550 4.000 122.030 4.280 ;
        RECT 123.150 4.000 127.550 4.280 ;
        RECT 128.670 4.000 132.150 4.280 ;
        RECT 133.270 4.000 136.750 4.280 ;
        RECT 137.870 4.000 141.350 4.280 ;
        RECT 142.470 4.000 145.950 4.280 ;
        RECT 147.070 4.000 150.550 4.280 ;
        RECT 151.670 4.000 155.150 4.280 ;
        RECT 156.270 4.000 160.670 4.280 ;
        RECT 161.790 4.000 165.270 4.280 ;
        RECT 166.390 4.000 169.870 4.280 ;
        RECT 170.990 4.000 174.470 4.280 ;
        RECT 175.590 4.000 179.070 4.280 ;
        RECT 180.190 4.000 183.670 4.280 ;
        RECT 184.790 4.000 189.190 4.280 ;
        RECT 190.310 4.000 193.790 4.280 ;
        RECT 194.910 4.000 198.390 4.280 ;
        RECT 199.510 4.000 202.990 4.280 ;
        RECT 204.110 4.000 207.590 4.280 ;
        RECT 208.710 4.000 212.190 4.280 ;
        RECT 213.310 4.000 216.790 4.280 ;
        RECT 217.910 4.000 222.310 4.280 ;
        RECT 223.430 4.000 226.910 4.280 ;
        RECT 228.030 4.000 231.510 4.280 ;
        RECT 232.630 4.000 236.110 4.280 ;
        RECT 237.230 4.000 240.710 4.280 ;
        RECT 241.830 4.000 245.310 4.280 ;
        RECT 246.430 4.000 250.830 4.280 ;
        RECT 251.950 4.000 255.430 4.280 ;
        RECT 256.550 4.000 260.030 4.280 ;
        RECT 261.150 4.000 264.630 4.280 ;
        RECT 265.750 4.000 269.230 4.280 ;
        RECT 270.350 4.000 273.830 4.280 ;
        RECT 274.950 4.000 278.430 4.280 ;
        RECT 279.550 4.000 283.950 4.280 ;
        RECT 285.070 4.000 288.550 4.280 ;
        RECT 289.670 4.000 293.150 4.280 ;
      LAYER met3 ;
        RECT 4.400 293.100 296.000 294.265 ;
        RECT 4.000 292.380 296.000 293.100 ;
        RECT 4.000 290.380 295.600 292.380 ;
        RECT 4.000 288.300 296.000 290.380 ;
        RECT 4.400 286.300 296.000 288.300 ;
        RECT 4.000 285.580 296.000 286.300 ;
        RECT 4.000 283.580 295.600 285.580 ;
        RECT 4.000 281.500 296.000 283.580 ;
        RECT 4.400 279.500 296.000 281.500 ;
        RECT 4.000 278.780 296.000 279.500 ;
        RECT 4.000 276.780 295.600 278.780 ;
        RECT 4.000 273.340 296.000 276.780 ;
        RECT 4.400 271.980 296.000 273.340 ;
        RECT 4.400 271.340 295.600 271.980 ;
        RECT 4.000 269.980 295.600 271.340 ;
        RECT 4.000 266.540 296.000 269.980 ;
        RECT 4.400 265.180 296.000 266.540 ;
        RECT 4.400 264.540 295.600 265.180 ;
        RECT 4.000 263.180 295.600 264.540 ;
        RECT 4.000 259.740 296.000 263.180 ;
        RECT 4.400 258.380 296.000 259.740 ;
        RECT 4.400 257.740 295.600 258.380 ;
        RECT 4.000 256.380 295.600 257.740 ;
        RECT 4.000 252.940 296.000 256.380 ;
        RECT 4.400 250.940 296.000 252.940 ;
        RECT 4.000 250.220 296.000 250.940 ;
        RECT 4.000 248.220 295.600 250.220 ;
        RECT 4.000 246.140 296.000 248.220 ;
        RECT 4.400 244.140 296.000 246.140 ;
        RECT 4.000 243.420 296.000 244.140 ;
        RECT 4.000 241.420 295.600 243.420 ;
        RECT 4.000 239.340 296.000 241.420 ;
        RECT 4.400 237.340 296.000 239.340 ;
        RECT 4.000 236.620 296.000 237.340 ;
        RECT 4.000 234.620 295.600 236.620 ;
        RECT 4.000 231.180 296.000 234.620 ;
        RECT 4.400 229.820 296.000 231.180 ;
        RECT 4.400 229.180 295.600 229.820 ;
        RECT 4.000 227.820 295.600 229.180 ;
        RECT 4.000 224.380 296.000 227.820 ;
        RECT 4.400 223.020 296.000 224.380 ;
        RECT 4.400 222.380 295.600 223.020 ;
        RECT 4.000 221.020 295.600 222.380 ;
        RECT 4.000 217.580 296.000 221.020 ;
        RECT 4.400 216.220 296.000 217.580 ;
        RECT 4.400 215.580 295.600 216.220 ;
        RECT 4.000 214.220 295.600 215.580 ;
        RECT 4.000 210.780 296.000 214.220 ;
        RECT 4.400 209.420 296.000 210.780 ;
        RECT 4.400 208.780 295.600 209.420 ;
        RECT 4.000 207.420 295.600 208.780 ;
        RECT 4.000 203.980 296.000 207.420 ;
        RECT 4.400 201.980 296.000 203.980 ;
        RECT 4.000 201.260 296.000 201.980 ;
        RECT 4.000 199.260 295.600 201.260 ;
        RECT 4.000 197.180 296.000 199.260 ;
        RECT 4.400 195.180 296.000 197.180 ;
        RECT 4.000 194.460 296.000 195.180 ;
        RECT 4.000 192.460 295.600 194.460 ;
        RECT 4.000 190.380 296.000 192.460 ;
        RECT 4.400 188.380 296.000 190.380 ;
        RECT 4.000 187.660 296.000 188.380 ;
        RECT 4.000 185.660 295.600 187.660 ;
        RECT 4.000 182.220 296.000 185.660 ;
        RECT 4.400 180.860 296.000 182.220 ;
        RECT 4.400 180.220 295.600 180.860 ;
        RECT 4.000 178.860 295.600 180.220 ;
        RECT 4.000 175.420 296.000 178.860 ;
        RECT 4.400 174.060 296.000 175.420 ;
        RECT 4.400 173.420 295.600 174.060 ;
        RECT 4.000 172.060 295.600 173.420 ;
        RECT 4.000 168.620 296.000 172.060 ;
        RECT 4.400 167.260 296.000 168.620 ;
        RECT 4.400 166.620 295.600 167.260 ;
        RECT 4.000 165.260 295.600 166.620 ;
        RECT 4.000 161.820 296.000 165.260 ;
        RECT 4.400 159.820 296.000 161.820 ;
        RECT 4.000 159.100 296.000 159.820 ;
        RECT 4.000 157.100 295.600 159.100 ;
        RECT 4.000 155.020 296.000 157.100 ;
        RECT 4.400 153.020 296.000 155.020 ;
        RECT 4.000 152.300 296.000 153.020 ;
        RECT 4.000 150.300 295.600 152.300 ;
        RECT 4.000 148.220 296.000 150.300 ;
        RECT 4.400 146.220 296.000 148.220 ;
        RECT 4.000 145.500 296.000 146.220 ;
        RECT 4.000 143.500 295.600 145.500 ;
        RECT 4.000 141.420 296.000 143.500 ;
        RECT 4.400 139.420 296.000 141.420 ;
        RECT 4.000 138.700 296.000 139.420 ;
        RECT 4.000 136.700 295.600 138.700 ;
        RECT 4.000 133.260 296.000 136.700 ;
        RECT 4.400 131.900 296.000 133.260 ;
        RECT 4.400 131.260 295.600 131.900 ;
        RECT 4.000 129.900 295.600 131.260 ;
        RECT 4.000 126.460 296.000 129.900 ;
        RECT 4.400 125.100 296.000 126.460 ;
        RECT 4.400 124.460 295.600 125.100 ;
        RECT 4.000 123.100 295.600 124.460 ;
        RECT 4.000 119.660 296.000 123.100 ;
        RECT 4.400 118.300 296.000 119.660 ;
        RECT 4.400 117.660 295.600 118.300 ;
        RECT 4.000 116.300 295.600 117.660 ;
        RECT 4.000 112.860 296.000 116.300 ;
        RECT 4.400 110.860 296.000 112.860 ;
        RECT 4.000 110.140 296.000 110.860 ;
        RECT 4.000 108.140 295.600 110.140 ;
        RECT 4.000 106.060 296.000 108.140 ;
        RECT 4.400 104.060 296.000 106.060 ;
        RECT 4.000 103.340 296.000 104.060 ;
        RECT 4.000 101.340 295.600 103.340 ;
        RECT 4.000 99.260 296.000 101.340 ;
        RECT 4.400 97.260 296.000 99.260 ;
        RECT 4.000 96.540 296.000 97.260 ;
        RECT 4.000 94.540 295.600 96.540 ;
        RECT 4.000 91.100 296.000 94.540 ;
        RECT 4.400 89.740 296.000 91.100 ;
        RECT 4.400 89.100 295.600 89.740 ;
        RECT 4.000 87.740 295.600 89.100 ;
        RECT 4.000 84.300 296.000 87.740 ;
        RECT 4.400 82.940 296.000 84.300 ;
        RECT 4.400 82.300 295.600 82.940 ;
        RECT 4.000 80.940 295.600 82.300 ;
        RECT 4.000 77.500 296.000 80.940 ;
        RECT 4.400 76.140 296.000 77.500 ;
        RECT 4.400 75.500 295.600 76.140 ;
        RECT 4.000 74.140 295.600 75.500 ;
        RECT 4.000 70.700 296.000 74.140 ;
        RECT 4.400 69.340 296.000 70.700 ;
        RECT 4.400 68.700 295.600 69.340 ;
        RECT 4.000 67.340 295.600 68.700 ;
        RECT 4.000 63.900 296.000 67.340 ;
        RECT 4.400 61.900 296.000 63.900 ;
        RECT 4.000 61.180 296.000 61.900 ;
        RECT 4.000 59.180 295.600 61.180 ;
        RECT 4.000 57.100 296.000 59.180 ;
        RECT 4.400 55.100 296.000 57.100 ;
        RECT 4.000 54.380 296.000 55.100 ;
        RECT 4.000 52.380 295.600 54.380 ;
        RECT 4.000 50.300 296.000 52.380 ;
        RECT 4.400 48.300 296.000 50.300 ;
        RECT 4.000 47.580 296.000 48.300 ;
        RECT 4.000 45.580 295.600 47.580 ;
        RECT 4.000 42.140 296.000 45.580 ;
        RECT 4.400 40.780 296.000 42.140 ;
        RECT 4.400 40.140 295.600 40.780 ;
        RECT 4.000 38.780 295.600 40.140 ;
        RECT 4.000 35.340 296.000 38.780 ;
        RECT 4.400 33.980 296.000 35.340 ;
        RECT 4.400 33.340 295.600 33.980 ;
        RECT 4.000 31.980 295.600 33.340 ;
        RECT 4.000 28.540 296.000 31.980 ;
        RECT 4.400 27.180 296.000 28.540 ;
        RECT 4.400 26.540 295.600 27.180 ;
        RECT 4.000 25.180 295.600 26.540 ;
        RECT 4.000 21.740 296.000 25.180 ;
        RECT 4.400 19.740 296.000 21.740 ;
        RECT 4.000 19.020 296.000 19.740 ;
        RECT 4.000 17.020 295.600 19.020 ;
        RECT 4.000 14.940 296.000 17.020 ;
        RECT 4.400 12.940 296.000 14.940 ;
        RECT 4.000 12.220 296.000 12.940 ;
        RECT 4.000 10.715 295.600 12.220 ;
  END
END wrapped_asic_watch
END LIBRARY

