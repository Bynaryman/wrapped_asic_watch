VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO wrapped_asic_watch
  CLASS BLOCK ;
  FOREIGN wrapped_asic_watch ;
  ORIGIN 0.000 0.000 ;
  SIZE 100.000 BY 220.000 ;
  PIN active
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 165.660 4.000 166.860 ;
    END
  END active
  PIN io_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 39.510 0.000 40.070 4.000 ;
    END
  END io_in[0]
  PIN io_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 43.190 216.000 43.750 220.000 ;
    END
  END io_in[10]
  PIN io_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 179.260 4.000 180.460 ;
    END
  END io_in[11]
  PIN io_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 96.000 191.500 100.000 192.700 ;
    END
  END io_in[12]
  PIN io_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 60.670 0.000 61.230 4.000 ;
    END
  END io_in[13]
  PIN io_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 20.190 216.000 20.750 220.000 ;
    END
  END io_in[14]
  PIN io_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 96.000 198.300 100.000 199.500 ;
    END
  END io_in[15]
  PIN io_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 96.000 55.500 100.000 56.700 ;
    END
  END io_in[16]
  PIN io_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 218.700 4.000 219.900 ;
    END
  END io_in[17]
  PIN io_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3.630 216.000 4.190 220.000 ;
    END
  END io_in[18]
  PIN io_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 96.000 14.700 100.000 15.900 ;
    END
  END io_in[19]
  PIN io_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 58.220 4.000 59.420 ;
    END
  END io_in[1]
  PIN io_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 103.100 4.000 104.300 ;
    END
  END io_in[20]
  PIN io_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 69.100 4.000 70.300 ;
    END
  END io_in[21]
  PIN io_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 96.000 97.660 100.000 98.860 ;
    END
  END io_in[22]
  PIN io_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 214.620 4.000 215.820 ;
    END
  END io_in[23]
  PIN io_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 203.740 4.000 204.940 ;
    END
  END io_in[24]
  PIN io_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 95.630 0.000 96.190 4.000 ;
    END
  END io_in[25]
  PIN io_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 93.790 0.000 94.350 4.000 ;
    END
  END io_in[26]
  PIN io_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 96.000 79.980 100.000 81.180 ;
    END
  END io_in[27]
  PIN io_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 84.590 0.000 85.150 4.000 ;
    END
  END io_in[28]
  PIN io_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 99.310 216.000 99.870 220.000 ;
    END
  END io_in[29]
  PIN io_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 42.270 0.000 42.830 4.000 ;
    END
  END io_in[2]
  PIN io_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 96.000 111.260 100.000 112.460 ;
    END
  END io_in[30]
  PIN io_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 158.860 4.000 160.060 ;
    END
  END io_in[31]
  PIN io_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 79.070 0.000 79.630 4.000 ;
    END
  END io_in[32]
  PIN io_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 93.580 4.000 94.780 ;
    END
  END io_in[33]
  PIN io_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 68.950 216.000 69.510 220.000 ;
    END
  END io_in[34]
  PIN io_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 83.670 216.000 84.230 220.000 ;
    END
  END io_in[35]
  PIN io_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 96.000 153.420 100.000 154.620 ;
    END
  END io_in[36]
  PIN io_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 85.510 216.000 86.070 220.000 ;
    END
  END io_in[37]
  PIN io_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 45.950 216.000 46.510 220.000 ;
    END
  END io_in[3]
  PIN io_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 96.000 149.340 100.000 150.540 ;
    END
  END io_in[4]
  PIN io_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 96.000 211.900 100.000 213.100 ;
    END
  END io_in[5]
  PIN io_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 109.900 4.000 111.100 ;
    END
  END io_in[6]
  PIN io_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 75.900 4.000 77.100 ;
    END
  END io_in[7]
  PIN io_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 96.000 160.220 100.000 161.420 ;
    END
  END io_in[8]
  PIN io_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 210.540 4.000 211.740 ;
    END
  END io_in[9]
  PIN io_oeb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 68.030 0.000 68.590 4.000 ;
    END
  END io_oeb[0]
  PIN io_oeb[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 62.300 4.000 63.500 ;
    END
  END io_oeb[10]
  PIN io_oeb[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 96.000 142.540 100.000 143.740 ;
    END
  END io_oeb[11]
  PIN io_oeb[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 96.000 93.580 100.000 94.780 ;
    END
  END io_oeb[12]
  PIN io_oeb[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 96.000 90.860 100.000 92.060 ;
    END
  END io_oeb[13]
  PIN io_oeb[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 16.060 4.000 17.260 ;
    END
  END io_oeb[14]
  PIN io_oeb[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 8.230 216.000 8.790 220.000 ;
    END
  END io_oeb[15]
  PIN io_oeb[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 96.000 48.700 100.000 49.900 ;
    END
  END io_oeb[16]
  PIN io_oeb[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 34.910 0.000 35.470 4.000 ;
    END
  END io_oeb[17]
  PIN io_oeb[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 64.350 216.000 64.910 220.000 ;
    END
  END io_oeb[18]
  PIN io_oeb[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 10.070 216.000 10.630 220.000 ;
    END
  END io_oeb[19]
  PIN io_oeb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 96.000 -0.260 100.000 0.940 ;
    END
  END io_oeb[1]
  PIN io_oeb[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 96.000 118.060 100.000 119.260 ;
    END
  END io_oeb[20]
  PIN io_oeb[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 187.420 4.000 188.620 ;
    END
  END io_oeb[21]
  PIN io_oeb[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 13.750 0.000 14.310 4.000 ;
    END
  END io_oeb[22]
  PIN io_oeb[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 35.830 216.000 36.390 220.000 ;
    END
  END io_oeb[23]
  PIN io_oeb[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 38.590 216.000 39.150 220.000 ;
    END
  END io_oeb[24]
  PIN io_oeb[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 96.000 31.020 100.000 32.220 ;
    END
  END io_oeb[25]
  PIN io_oeb[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 96.000 180.620 100.000 181.820 ;
    END
  END io_oeb[26]
  PIN io_oeb[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 47.790 216.000 48.350 220.000 ;
    END
  END io_oeb[27]
  PIN io_oeb[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 96.000 10.620 100.000 11.820 ;
    END
  END io_oeb[28]
  PIN io_oeb[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 96.000 156.140 100.000 157.340 ;
    END
  END io_oeb[29]
  PIN io_oeb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 78.150 216.000 78.710 220.000 ;
    END
  END io_oeb[2]
  PIN io_oeb[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 190.140 4.000 191.340 ;
    END
  END io_oeb[30]
  PIN io_oeb[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 96.000 7.900 100.000 9.100 ;
    END
  END io_oeb[31]
  PIN io_oeb[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 89.500 4.000 90.700 ;
    END
  END io_oeb[32]
  PIN io_oeb[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 96.000 35.100 100.000 36.300 ;
    END
  END io_oeb[33]
  PIN io_oeb[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.870 216.000 1.430 220.000 ;
    END
  END io_oeb[34]
  PIN io_oeb[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 78.620 4.000 79.820 ;
    END
  END io_oeb[35]
  PIN io_oeb[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 40.540 4.000 41.740 ;
    END
  END io_oeb[36]
  PIN io_oeb[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 65.020 4.000 66.220 ;
    END
  END io_oeb[37]
  PIN io_oeb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 65.270 0.000 65.830 4.000 ;
    END
  END io_oeb[3]
  PIN io_oeb[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 96.000 41.900 100.000 43.100 ;
    END
  END io_oeb[4]
  PIN io_oeb[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 116.700 4.000 117.900 ;
    END
  END io_oeb[5]
  PIN io_oeb[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 96.000 104.460 100.000 105.660 ;
    END
  END io_oeb[6]
  PIN io_oeb[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 5.470 216.000 6.030 220.000 ;
    END
  END io_oeb[7]
  PIN io_oeb[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 10.990 0.000 11.550 4.000 ;
    END
  END io_oeb[8]
  PIN io_oeb[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 27.550 0.000 28.110 4.000 ;
    END
  END io_oeb[9]
  PIN io_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 96.000 209.180 100.000 210.380 ;
    END
  END io_out[0]
  PIN io_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 96.000 139.820 100.000 141.020 ;
    END
  END io_out[10]
  PIN io_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 9.260 4.000 10.460 ;
    END
  END io_out[11]
  PIN io_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 26.940 4.000 28.140 ;
    END
  END io_out[12]
  PIN io_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 96.000 3.820 100.000 5.020 ;
    END
  END io_out[13]
  PIN io_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 96.000 184.700 100.000 185.900 ;
    END
  END io_out[14]
  PIN io_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 147.980 4.000 149.180 ;
    END
  END io_out[15]
  PIN io_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 96.000 135.740 100.000 136.940 ;
    END
  END io_out[16]
  PIN io_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 90.110 216.000 90.670 220.000 ;
    END
  END io_out[17]
  PIN io_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 96.000 28.300 100.000 29.500 ;
    END
  END io_out[18]
  PIN io_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 85.420 4.000 86.620 ;
    END
  END io_out[19]
  PIN io_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 56.990 216.000 57.550 220.000 ;
    END
  END io_out[1]
  PIN io_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 76.310 216.000 76.870 220.000 ;
    END
  END io_out[20]
  PIN io_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 145.260 4.000 146.460 ;
    END
  END io_out[21]
  PIN io_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 81.830 0.000 82.390 4.000 ;
    END
  END io_out[22]
  PIN io_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 96.000 122.140 100.000 123.340 ;
    END
  END io_out[23]
  PIN io_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 69.870 0.000 70.430 4.000 ;
    END
  END io_out[24]
  PIN io_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 67.110 216.000 67.670 220.000 ;
    END
  END io_out[25]
  PIN io_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 20.140 4.000 21.340 ;
    END
  END io_out[26]
  PIN io_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 71.710 216.000 72.270 220.000 ;
    END
  END io_out[27]
  PIN io_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 44.110 0.000 44.670 4.000 ;
    END
  END io_out[28]
  PIN io_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 96.000 45.980 100.000 47.180 ;
    END
  END io_out[29]
  PIN io_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 18.350 0.000 18.910 4.000 ;
    END
  END io_out[2]
  PIN io_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 22.860 4.000 24.060 ;
    END
  END io_out[30]
  PIN io_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 51.420 4.000 52.620 ;
    END
  END io_out[31]
  PIN io_out[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 169.740 4.000 170.940 ;
    END
  END io_out[32]
  PIN io_out[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 96.000 66.380 100.000 67.580 ;
    END
  END io_out[33]
  PIN io_out[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 96.000 187.420 100.000 188.620 ;
    END
  END io_out[34]
  PIN io_out[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 96.000 177.900 100.000 179.100 ;
    END
  END io_out[35]
  PIN io_out[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 12.830 216.000 13.390 220.000 ;
    END
  END io_out[36]
  PIN io_out[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 96.000 202.380 100.000 203.580 ;
    END
  END io_out[37]
  PIN io_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 156.140 4.000 157.340 ;
    END
  END io_out[3]
  PIN io_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 96.000 146.620 100.000 147.820 ;
    END
  END io_out[4]
  PIN io_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 31.230 216.000 31.790 220.000 ;
    END
  END io_out[5]
  PIN io_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 94.710 216.000 95.270 220.000 ;
    END
  END io_out[6]
  PIN io_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 71.820 4.000 73.020 ;
    END
  END io_out[7]
  PIN io_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 48.710 0.000 49.270 4.000 ;
    END
  END io_out[8]
  PIN io_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 54.140 4.000 55.340 ;
    END
  END io_out[9]
  PIN la1_data_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 96.000 70.460 100.000 71.660 ;
    END
  END la1_data_in[0]
  PIN la1_data_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 56.070 0.000 56.630 4.000 ;
    END
  END la1_data_in[10]
  PIN la1_data_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 96.000 62.300 100.000 63.500 ;
    END
  END la1_data_in[11]
  PIN la1_data_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 134.380 4.000 135.580 ;
    END
  END la1_data_in[12]
  PIN la1_data_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 86.430 0.000 86.990 4.000 ;
    END
  END la1_data_in[13]
  PIN la1_data_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 47.340 4.000 48.540 ;
    END
  END la1_data_in[14]
  PIN la1_data_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 14.670 216.000 15.230 220.000 ;
    END
  END la1_data_in[15]
  PIN la1_data_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 52.390 216.000 52.950 220.000 ;
    END
  END la1_data_in[16]
  PIN la1_data_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 33.990 216.000 34.550 220.000 ;
    END
  END la1_data_in[17]
  PIN la1_data_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 96.000 17.420 100.000 18.620 ;
    END
  END la1_data_in[18]
  PIN la1_data_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 17.430 216.000 17.990 220.000 ;
    END
  END la1_data_in[19]
  PIN la1_data_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 51.470 0.000 52.030 4.000 ;
    END
  END la1_data_in[1]
  PIN la1_data_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 131.660 4.000 132.860 ;
    END
  END la1_data_in[20]
  PIN la1_data_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 97.470 216.000 98.030 220.000 ;
    END
  END la1_data_in[21]
  PIN la1_data_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 96.000 73.180 100.000 74.380 ;
    END
  END la1_data_in[22]
  PIN la1_data_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2.460 4.000 3.660 ;
    END
  END la1_data_in[23]
  PIN la1_data_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 36.750 0.000 37.310 4.000 ;
    END
  END la1_data_in[24]
  PIN la1_data_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 138.460 4.000 139.660 ;
    END
  END la1_data_in[25]
  PIN la1_data_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 96.000 52.780 100.000 53.980 ;
    END
  END la1_data_in[26]
  PIN la1_data_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 74.470 0.000 75.030 4.000 ;
    END
  END la1_data_in[27]
  PIN la1_data_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 120.780 4.000 121.980 ;
    END
  END la1_data_in[28]
  PIN la1_data_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 183.340 4.000 184.540 ;
    END
  END la1_data_in[29]
  PIN la1_data_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 30.310 0.000 30.870 4.000 ;
    END
  END la1_data_in[2]
  PIN la1_data_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 4.550 0.000 5.110 4.000 ;
    END
  END la1_data_in[30]
  PIN la1_data_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 98.390 0.000 98.950 4.000 ;
    END
  END la1_data_in[31]
  PIN la1_data_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 113.980 4.000 115.180 ;
    END
  END la1_data_in[3]
  PIN la1_data_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 80.910 216.000 81.470 220.000 ;
    END
  END la1_data_in[4]
  PIN la1_data_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 96.000 128.940 100.000 130.140 ;
    END
  END la1_data_in[5]
  PIN la1_data_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 22.030 216.000 22.590 220.000 ;
    END
  END la1_data_in[6]
  PIN la1_data_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 82.700 4.000 83.900 ;
    END
  END la1_data_in[7]
  PIN la1_data_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 24.790 216.000 25.350 220.000 ;
    END
  END la1_data_in[8]
  PIN la1_data_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 124.860 4.000 126.060 ;
    END
  END la1_data_in[9]
  PIN la1_data_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 21.110 0.000 21.670 4.000 ;
    END
  END la1_data_out[0]
  PIN la1_data_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 96.000 84.060 100.000 85.260 ;
    END
  END la1_data_out[10]
  PIN la1_data_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 57.910 0.000 58.470 4.000 ;
    END
  END la1_data_out[11]
  PIN la1_data_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 96.000 205.100 100.000 206.300 ;
    END
  END la1_data_out[12]
  PIN la1_data_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 196.940 4.000 198.140 ;
    END
  END la1_data_out[13]
  PIN la1_data_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 41.350 216.000 41.910 220.000 ;
    END
  END la1_data_out[14]
  PIN la1_data_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 6.540 4.000 7.740 ;
    END
  END la1_data_out[15]
  PIN la1_data_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 96.000 101.740 100.000 102.940 ;
    END
  END la1_data_out[16]
  PIN la1_data_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 96.000 171.100 100.000 172.300 ;
    END
  END la1_data_out[17]
  PIN la1_data_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 201.020 4.000 202.220 ;
    END
  END la1_data_out[18]
  PIN la1_data_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 96.000 133.020 100.000 134.220 ;
    END
  END la1_data_out[19]
  PIN la1_data_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 162.940 4.000 164.140 ;
    END
  END la1_data_out[1]
  PIN la1_data_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 37.820 4.000 39.020 ;
    END
  END la1_data_out[20]
  PIN la1_data_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 96.000 195.580 100.000 196.780 ;
    END
  END la1_data_out[21]
  PIN la1_data_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 50.550 216.000 51.110 220.000 ;
    END
  END la1_data_out[22]
  PIN la1_data_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 32.150 0.000 32.710 4.000 ;
    END
  END la1_data_out[23]
  PIN la1_data_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 96.000 108.540 100.000 109.740 ;
    END
  END la1_data_out[24]
  PIN la1_data_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 13.340 4.000 14.540 ;
    END
  END la1_data_out[25]
  PIN la1_data_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 96.000 59.580 100.000 60.780 ;
    END
  END la1_data_out[26]
  PIN la1_data_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 172.460 4.000 173.660 ;
    END
  END la1_data_out[27]
  PIN la1_data_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 96.000 21.500 100.000 22.700 ;
    END
  END la1_data_out[28]
  PIN la1_data_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 15.590 0.000 16.150 4.000 ;
    END
  END la1_data_out[29]
  PIN la1_data_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 53.310 0.000 53.870 4.000 ;
    END
  END la1_data_out[2]
  PIN la1_data_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 96.000 86.780 100.000 87.980 ;
    END
  END la1_data_out[30]
  PIN la1_data_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 96.000 215.980 100.000 217.180 ;
    END
  END la1_data_out[31]
  PIN la1_data_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 33.740 4.000 34.940 ;
    END
  END la1_data_out[3]
  PIN la1_data_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 96.000 24.220 100.000 25.420 ;
    END
  END la1_data_out[4]
  PIN la1_data_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 9.150 0.000 9.710 4.000 ;
    END
  END la1_data_out[5]
  PIN la1_data_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 96.000 115.340 100.000 116.540 ;
    END
  END la1_data_out[6]
  PIN la1_data_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1.790 0.000 2.350 4.000 ;
    END
  END la1_data_out[7]
  PIN la1_data_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 96.000 173.820 100.000 175.020 ;
    END
  END la1_data_out[8]
  PIN la1_data_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 92.870 216.000 93.430 220.000 ;
    END
  END la1_data_out[9]
  PIN la1_oenb[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 96.000 39.180 100.000 40.380 ;
    END
  END la1_oenb[0]
  PIN la1_oenb[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 88.270 216.000 88.830 220.000 ;
    END
  END la1_oenb[10]
  PIN la1_oenb[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 100.380 4.000 101.580 ;
    END
  END la1_oenb[11]
  PIN la1_oenb[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 107.180 4.000 108.380 ;
    END
  END la1_oenb[12]
  PIN la1_oenb[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 77.230 0.000 77.790 4.000 ;
    END
  END la1_oenb[13]
  PIN la1_oenb[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT -0.050 0.000 0.510 4.000 ;
    END
  END la1_oenb[14]
  PIN la1_oenb[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 91.030 0.000 91.590 4.000 ;
    END
  END la1_oenb[15]
  PIN la1_oenb[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 127.580 4.000 128.780 ;
    END
  END la1_oenb[16]
  PIN la1_oenb[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 194.220 4.000 195.420 ;
    END
  END la1_oenb[17]
  PIN la1_oenb[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 29.390 216.000 29.950 220.000 ;
    END
  END la1_oenb[18]
  PIN la1_oenb[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 96.300 4.000 97.500 ;
    END
  END la1_oenb[19]
  PIN la1_oenb[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 22.950 0.000 23.510 4.000 ;
    END
  END la1_oenb[1]
  PIN la1_oenb[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 6.390 0.000 6.950 4.000 ;
    END
  END la1_oenb[20]
  PIN la1_oenb[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 55.150 216.000 55.710 220.000 ;
    END
  END la1_oenb[21]
  PIN la1_oenb[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 26.630 216.000 27.190 220.000 ;
    END
  END la1_oenb[22]
  PIN la1_oenb[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 63.430 0.000 63.990 4.000 ;
    END
  END la1_oenb[23]
  PIN la1_oenb[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 73.550 216.000 74.110 220.000 ;
    END
  END la1_oenb[24]
  PIN la1_oenb[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 96.000 77.260 100.000 78.460 ;
    END
  END la1_oenb[25]
  PIN la1_oenb[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 141.180 4.000 142.380 ;
    END
  END la1_oenb[26]
  PIN la1_oenb[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 96.000 167.020 100.000 168.220 ;
    END
  END la1_oenb[27]
  PIN la1_oenb[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 25.710 0.000 26.270 4.000 ;
    END
  END la1_oenb[28]
  PIN la1_oenb[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 46.870 0.000 47.430 4.000 ;
    END
  END la1_oenb[29]
  PIN la1_oenb[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 31.020 4.000 32.220 ;
    END
  END la1_oenb[2]
  PIN la1_oenb[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 96.000 164.300 100.000 165.500 ;
    END
  END la1_oenb[30]
  PIN la1_oenb[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 72.630 0.000 73.190 4.000 ;
    END
  END la1_oenb[31]
  PIN la1_oenb[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 62.510 216.000 63.070 220.000 ;
    END
  END la1_oenb[3]
  PIN la1_oenb[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 59.750 216.000 60.310 220.000 ;
    END
  END la1_oenb[4]
  PIN la1_oenb[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 176.540 4.000 177.740 ;
    END
  END la1_oenb[5]
  PIN la1_oenb[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 207.820 4.000 209.020 ;
    END
  END la1_oenb[6]
  PIN la1_oenb[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 89.190 0.000 89.750 4.000 ;
    END
  END la1_oenb[7]
  PIN la1_oenb[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 44.620 4.000 45.820 ;
    END
  END la1_oenb[8]
  PIN la1_oenb[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 152.060 4.000 153.260 ;
    END
  END la1_oenb[9]
  PIN vccd1
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 19.545 10.640 21.145 206.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 49.195 10.640 50.795 206.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 78.850 10.640 80.450 206.960 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 34.370 10.640 35.970 206.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 64.025 10.640 65.625 206.960 ;
    END
  END vssd1
  PIN wb_clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 96.000 124.860 100.000 126.060 ;
    END
  END wb_clk_i
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 95.075 206.805 ;
      LAYER met1 ;
        RECT 0.990 10.640 95.150 206.960 ;
      LAYER met2 ;
        RECT 1.710 215.720 3.350 216.765 ;
        RECT 4.470 215.720 5.190 216.765 ;
        RECT 6.310 215.720 7.950 216.765 ;
        RECT 9.070 215.720 9.790 216.765 ;
        RECT 10.910 215.720 12.550 216.765 ;
        RECT 13.670 215.720 14.390 216.765 ;
        RECT 15.510 215.720 17.150 216.765 ;
        RECT 18.270 215.720 19.910 216.765 ;
        RECT 21.030 215.720 21.750 216.765 ;
        RECT 22.870 215.720 24.510 216.765 ;
        RECT 25.630 215.720 26.350 216.765 ;
        RECT 27.470 215.720 29.110 216.765 ;
        RECT 30.230 215.720 30.950 216.765 ;
        RECT 32.070 215.720 33.710 216.765 ;
        RECT 34.830 215.720 35.550 216.765 ;
        RECT 36.670 215.720 38.310 216.765 ;
        RECT 39.430 215.720 41.070 216.765 ;
        RECT 42.190 215.720 42.910 216.765 ;
        RECT 44.030 215.720 45.670 216.765 ;
        RECT 46.790 215.720 47.510 216.765 ;
        RECT 48.630 215.720 50.270 216.765 ;
        RECT 51.390 215.720 52.110 216.765 ;
        RECT 53.230 215.720 54.870 216.765 ;
        RECT 55.990 215.720 56.710 216.765 ;
        RECT 57.830 215.720 59.470 216.765 ;
        RECT 60.590 215.720 62.230 216.765 ;
        RECT 63.350 215.720 64.070 216.765 ;
        RECT 65.190 215.720 66.830 216.765 ;
        RECT 67.950 215.720 68.670 216.765 ;
        RECT 69.790 215.720 71.430 216.765 ;
        RECT 72.550 215.720 73.270 216.765 ;
        RECT 74.390 215.720 76.030 216.765 ;
        RECT 77.150 215.720 77.870 216.765 ;
        RECT 78.990 215.720 80.630 216.765 ;
        RECT 81.750 215.720 83.390 216.765 ;
        RECT 84.510 215.720 85.230 216.765 ;
        RECT 86.350 215.720 87.990 216.765 ;
        RECT 89.110 215.720 89.830 216.765 ;
        RECT 90.950 215.720 92.590 216.765 ;
        RECT 93.710 215.720 94.430 216.765 ;
        RECT 1.020 4.280 95.120 215.720 ;
        RECT 1.020 0.155 1.510 4.280 ;
        RECT 2.630 0.155 4.270 4.280 ;
        RECT 5.390 0.155 6.110 4.280 ;
        RECT 7.230 0.155 8.870 4.280 ;
        RECT 9.990 0.155 10.710 4.280 ;
        RECT 11.830 0.155 13.470 4.280 ;
        RECT 14.590 0.155 15.310 4.280 ;
        RECT 16.430 0.155 18.070 4.280 ;
        RECT 19.190 0.155 20.830 4.280 ;
        RECT 21.950 0.155 22.670 4.280 ;
        RECT 23.790 0.155 25.430 4.280 ;
        RECT 26.550 0.155 27.270 4.280 ;
        RECT 28.390 0.155 30.030 4.280 ;
        RECT 31.150 0.155 31.870 4.280 ;
        RECT 32.990 0.155 34.630 4.280 ;
        RECT 35.750 0.155 36.470 4.280 ;
        RECT 37.590 0.155 39.230 4.280 ;
        RECT 40.350 0.155 41.990 4.280 ;
        RECT 43.110 0.155 43.830 4.280 ;
        RECT 44.950 0.155 46.590 4.280 ;
        RECT 47.710 0.155 48.430 4.280 ;
        RECT 49.550 0.155 51.190 4.280 ;
        RECT 52.310 0.155 53.030 4.280 ;
        RECT 54.150 0.155 55.790 4.280 ;
        RECT 56.910 0.155 57.630 4.280 ;
        RECT 58.750 0.155 60.390 4.280 ;
        RECT 61.510 0.155 63.150 4.280 ;
        RECT 64.270 0.155 64.990 4.280 ;
        RECT 66.110 0.155 67.750 4.280 ;
        RECT 68.870 0.155 69.590 4.280 ;
        RECT 70.710 0.155 72.350 4.280 ;
        RECT 73.470 0.155 74.190 4.280 ;
        RECT 75.310 0.155 76.950 4.280 ;
        RECT 78.070 0.155 78.790 4.280 ;
        RECT 79.910 0.155 81.550 4.280 ;
        RECT 82.670 0.155 84.310 4.280 ;
        RECT 85.430 0.155 86.150 4.280 ;
        RECT 87.270 0.155 88.910 4.280 ;
        RECT 90.030 0.155 90.750 4.280 ;
        RECT 91.870 0.155 93.510 4.280 ;
        RECT 94.630 0.155 95.120 4.280 ;
      LAYER met3 ;
        RECT 4.000 216.220 95.600 216.745 ;
        RECT 4.400 215.580 95.600 216.220 ;
        RECT 4.400 214.220 96.000 215.580 ;
        RECT 4.000 213.500 96.000 214.220 ;
        RECT 4.000 212.140 95.600 213.500 ;
        RECT 4.400 211.500 95.600 212.140 ;
        RECT 4.400 210.780 96.000 211.500 ;
        RECT 4.400 210.140 95.600 210.780 ;
        RECT 4.000 209.420 95.600 210.140 ;
        RECT 4.400 208.780 95.600 209.420 ;
        RECT 4.400 207.420 96.000 208.780 ;
        RECT 4.000 206.700 96.000 207.420 ;
        RECT 4.000 205.340 95.600 206.700 ;
        RECT 4.400 204.700 95.600 205.340 ;
        RECT 4.400 203.980 96.000 204.700 ;
        RECT 4.400 203.340 95.600 203.980 ;
        RECT 4.000 202.620 95.600 203.340 ;
        RECT 4.400 201.980 95.600 202.620 ;
        RECT 4.400 200.620 96.000 201.980 ;
        RECT 4.000 199.900 96.000 200.620 ;
        RECT 4.000 198.540 95.600 199.900 ;
        RECT 4.400 197.900 95.600 198.540 ;
        RECT 4.400 197.180 96.000 197.900 ;
        RECT 4.400 196.540 95.600 197.180 ;
        RECT 4.000 195.820 95.600 196.540 ;
        RECT 4.400 195.180 95.600 195.820 ;
        RECT 4.400 193.820 96.000 195.180 ;
        RECT 4.000 193.100 96.000 193.820 ;
        RECT 4.000 191.740 95.600 193.100 ;
        RECT 4.400 191.100 95.600 191.740 ;
        RECT 4.400 189.740 96.000 191.100 ;
        RECT 4.000 189.020 96.000 189.740 ;
        RECT 4.400 187.020 95.600 189.020 ;
        RECT 4.000 186.300 96.000 187.020 ;
        RECT 4.000 184.940 95.600 186.300 ;
        RECT 4.400 184.300 95.600 184.940 ;
        RECT 4.400 182.940 96.000 184.300 ;
        RECT 4.000 182.220 96.000 182.940 ;
        RECT 4.000 180.860 95.600 182.220 ;
        RECT 4.400 180.220 95.600 180.860 ;
        RECT 4.400 179.500 96.000 180.220 ;
        RECT 4.400 178.860 95.600 179.500 ;
        RECT 4.000 178.140 95.600 178.860 ;
        RECT 4.400 177.500 95.600 178.140 ;
        RECT 4.400 176.140 96.000 177.500 ;
        RECT 4.000 175.420 96.000 176.140 ;
        RECT 4.000 174.060 95.600 175.420 ;
        RECT 4.400 173.420 95.600 174.060 ;
        RECT 4.400 172.700 96.000 173.420 ;
        RECT 4.400 172.060 95.600 172.700 ;
        RECT 4.000 171.340 95.600 172.060 ;
        RECT 4.400 170.700 95.600 171.340 ;
        RECT 4.400 169.340 96.000 170.700 ;
        RECT 4.000 168.620 96.000 169.340 ;
        RECT 4.000 167.260 95.600 168.620 ;
        RECT 4.400 166.620 95.600 167.260 ;
        RECT 4.400 165.900 96.000 166.620 ;
        RECT 4.400 165.260 95.600 165.900 ;
        RECT 4.000 164.540 95.600 165.260 ;
        RECT 4.400 163.900 95.600 164.540 ;
        RECT 4.400 162.540 96.000 163.900 ;
        RECT 4.000 161.820 96.000 162.540 ;
        RECT 4.000 160.460 95.600 161.820 ;
        RECT 4.400 159.820 95.600 160.460 ;
        RECT 4.400 158.460 96.000 159.820 ;
        RECT 4.000 157.740 96.000 158.460 ;
        RECT 4.400 155.740 95.600 157.740 ;
        RECT 4.000 155.020 96.000 155.740 ;
        RECT 4.000 153.660 95.600 155.020 ;
        RECT 4.400 153.020 95.600 153.660 ;
        RECT 4.400 151.660 96.000 153.020 ;
        RECT 4.000 150.940 96.000 151.660 ;
        RECT 4.000 149.580 95.600 150.940 ;
        RECT 4.400 148.940 95.600 149.580 ;
        RECT 4.400 148.220 96.000 148.940 ;
        RECT 4.400 147.580 95.600 148.220 ;
        RECT 4.000 146.860 95.600 147.580 ;
        RECT 4.400 146.220 95.600 146.860 ;
        RECT 4.400 144.860 96.000 146.220 ;
        RECT 4.000 144.140 96.000 144.860 ;
        RECT 4.000 142.780 95.600 144.140 ;
        RECT 4.400 142.140 95.600 142.780 ;
        RECT 4.400 141.420 96.000 142.140 ;
        RECT 4.400 140.780 95.600 141.420 ;
        RECT 4.000 140.060 95.600 140.780 ;
        RECT 4.400 139.420 95.600 140.060 ;
        RECT 4.400 138.060 96.000 139.420 ;
        RECT 4.000 137.340 96.000 138.060 ;
        RECT 4.000 135.980 95.600 137.340 ;
        RECT 4.400 135.340 95.600 135.980 ;
        RECT 4.400 134.620 96.000 135.340 ;
        RECT 4.400 133.980 95.600 134.620 ;
        RECT 4.000 133.260 95.600 133.980 ;
        RECT 4.400 132.620 95.600 133.260 ;
        RECT 4.400 131.260 96.000 132.620 ;
        RECT 4.000 130.540 96.000 131.260 ;
        RECT 4.000 129.180 95.600 130.540 ;
        RECT 4.400 128.540 95.600 129.180 ;
        RECT 4.400 127.180 96.000 128.540 ;
        RECT 4.000 126.460 96.000 127.180 ;
        RECT 4.400 124.460 95.600 126.460 ;
        RECT 4.000 123.740 96.000 124.460 ;
        RECT 4.000 122.380 95.600 123.740 ;
        RECT 4.400 121.740 95.600 122.380 ;
        RECT 4.400 120.380 96.000 121.740 ;
        RECT 4.000 119.660 96.000 120.380 ;
        RECT 4.000 118.300 95.600 119.660 ;
        RECT 4.400 117.660 95.600 118.300 ;
        RECT 4.400 116.940 96.000 117.660 ;
        RECT 4.400 116.300 95.600 116.940 ;
        RECT 4.000 115.580 95.600 116.300 ;
        RECT 4.400 114.940 95.600 115.580 ;
        RECT 4.400 113.580 96.000 114.940 ;
        RECT 4.000 112.860 96.000 113.580 ;
        RECT 4.000 111.500 95.600 112.860 ;
        RECT 4.400 110.860 95.600 111.500 ;
        RECT 4.400 110.140 96.000 110.860 ;
        RECT 4.400 109.500 95.600 110.140 ;
        RECT 4.000 108.780 95.600 109.500 ;
        RECT 4.400 108.140 95.600 108.780 ;
        RECT 4.400 106.780 96.000 108.140 ;
        RECT 4.000 106.060 96.000 106.780 ;
        RECT 4.000 104.700 95.600 106.060 ;
        RECT 4.400 104.060 95.600 104.700 ;
        RECT 4.400 103.340 96.000 104.060 ;
        RECT 4.400 102.700 95.600 103.340 ;
        RECT 4.000 101.980 95.600 102.700 ;
        RECT 4.400 101.340 95.600 101.980 ;
        RECT 4.400 99.980 96.000 101.340 ;
        RECT 4.000 99.260 96.000 99.980 ;
        RECT 4.000 97.900 95.600 99.260 ;
        RECT 4.400 97.260 95.600 97.900 ;
        RECT 4.400 95.900 96.000 97.260 ;
        RECT 4.000 95.180 96.000 95.900 ;
        RECT 4.400 93.180 95.600 95.180 ;
        RECT 4.000 92.460 96.000 93.180 ;
        RECT 4.000 91.100 95.600 92.460 ;
        RECT 4.400 90.460 95.600 91.100 ;
        RECT 4.400 89.100 96.000 90.460 ;
        RECT 4.000 88.380 96.000 89.100 ;
        RECT 4.000 87.020 95.600 88.380 ;
        RECT 4.400 86.380 95.600 87.020 ;
        RECT 4.400 85.660 96.000 86.380 ;
        RECT 4.400 85.020 95.600 85.660 ;
        RECT 4.000 84.300 95.600 85.020 ;
        RECT 4.400 83.660 95.600 84.300 ;
        RECT 4.400 82.300 96.000 83.660 ;
        RECT 4.000 81.580 96.000 82.300 ;
        RECT 4.000 80.220 95.600 81.580 ;
        RECT 4.400 79.580 95.600 80.220 ;
        RECT 4.400 78.860 96.000 79.580 ;
        RECT 4.400 78.220 95.600 78.860 ;
        RECT 4.000 77.500 95.600 78.220 ;
        RECT 4.400 76.860 95.600 77.500 ;
        RECT 4.400 75.500 96.000 76.860 ;
        RECT 4.000 74.780 96.000 75.500 ;
        RECT 4.000 73.420 95.600 74.780 ;
        RECT 4.400 72.780 95.600 73.420 ;
        RECT 4.400 72.060 96.000 72.780 ;
        RECT 4.400 71.420 95.600 72.060 ;
        RECT 4.000 70.700 95.600 71.420 ;
        RECT 4.400 70.060 95.600 70.700 ;
        RECT 4.400 68.700 96.000 70.060 ;
        RECT 4.000 67.980 96.000 68.700 ;
        RECT 4.000 66.620 95.600 67.980 ;
        RECT 4.400 65.980 95.600 66.620 ;
        RECT 4.400 64.620 96.000 65.980 ;
        RECT 4.000 63.900 96.000 64.620 ;
        RECT 4.400 61.900 95.600 63.900 ;
        RECT 4.000 61.180 96.000 61.900 ;
        RECT 4.000 59.820 95.600 61.180 ;
        RECT 4.400 59.180 95.600 59.820 ;
        RECT 4.400 57.820 96.000 59.180 ;
        RECT 4.000 57.100 96.000 57.820 ;
        RECT 4.000 55.740 95.600 57.100 ;
        RECT 4.400 55.100 95.600 55.740 ;
        RECT 4.400 54.380 96.000 55.100 ;
        RECT 4.400 53.740 95.600 54.380 ;
        RECT 4.000 53.020 95.600 53.740 ;
        RECT 4.400 52.380 95.600 53.020 ;
        RECT 4.400 51.020 96.000 52.380 ;
        RECT 4.000 50.300 96.000 51.020 ;
        RECT 4.000 48.940 95.600 50.300 ;
        RECT 4.400 48.300 95.600 48.940 ;
        RECT 4.400 47.580 96.000 48.300 ;
        RECT 4.400 46.940 95.600 47.580 ;
        RECT 4.000 46.220 95.600 46.940 ;
        RECT 4.400 45.580 95.600 46.220 ;
        RECT 4.400 44.220 96.000 45.580 ;
        RECT 4.000 43.500 96.000 44.220 ;
        RECT 4.000 42.140 95.600 43.500 ;
        RECT 4.400 41.500 95.600 42.140 ;
        RECT 4.400 40.780 96.000 41.500 ;
        RECT 4.400 40.140 95.600 40.780 ;
        RECT 4.000 39.420 95.600 40.140 ;
        RECT 4.400 38.780 95.600 39.420 ;
        RECT 4.400 37.420 96.000 38.780 ;
        RECT 4.000 36.700 96.000 37.420 ;
        RECT 4.000 35.340 95.600 36.700 ;
        RECT 4.400 34.700 95.600 35.340 ;
        RECT 4.400 33.340 96.000 34.700 ;
        RECT 4.000 32.620 96.000 33.340 ;
        RECT 4.400 30.620 95.600 32.620 ;
        RECT 4.000 29.900 96.000 30.620 ;
        RECT 4.000 28.540 95.600 29.900 ;
        RECT 4.400 27.900 95.600 28.540 ;
        RECT 4.400 26.540 96.000 27.900 ;
        RECT 4.000 25.820 96.000 26.540 ;
        RECT 4.000 24.460 95.600 25.820 ;
        RECT 4.400 23.820 95.600 24.460 ;
        RECT 4.400 23.100 96.000 23.820 ;
        RECT 4.400 22.460 95.600 23.100 ;
        RECT 4.000 21.740 95.600 22.460 ;
        RECT 4.400 21.100 95.600 21.740 ;
        RECT 4.400 19.740 96.000 21.100 ;
        RECT 4.000 19.020 96.000 19.740 ;
        RECT 4.000 17.660 95.600 19.020 ;
        RECT 4.400 17.020 95.600 17.660 ;
        RECT 4.400 16.300 96.000 17.020 ;
        RECT 4.400 15.660 95.600 16.300 ;
        RECT 4.000 14.940 95.600 15.660 ;
        RECT 4.400 14.300 95.600 14.940 ;
        RECT 4.400 12.940 96.000 14.300 ;
        RECT 4.000 12.220 96.000 12.940 ;
        RECT 4.000 10.860 95.600 12.220 ;
        RECT 4.400 10.220 95.600 10.860 ;
        RECT 4.400 9.500 96.000 10.220 ;
        RECT 4.400 8.860 95.600 9.500 ;
        RECT 4.000 8.140 95.600 8.860 ;
        RECT 4.400 7.500 95.600 8.140 ;
        RECT 4.400 6.140 96.000 7.500 ;
        RECT 4.000 5.420 96.000 6.140 ;
        RECT 4.000 4.060 95.600 5.420 ;
        RECT 4.400 3.420 95.600 4.060 ;
        RECT 4.400 2.060 96.000 3.420 ;
        RECT 4.000 1.340 96.000 2.060 ;
        RECT 4.000 0.175 95.600 1.340 ;
  END
END wrapped_asic_watch
END LIBRARY

